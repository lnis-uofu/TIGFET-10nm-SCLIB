* sclib_tigfet10_hpnw8_tt_0p70v_25c.sp
.subckt TIGFET_HPNW8 D PGD CG PGS S
xgate (D PGD CG PGS S) TIGFET nw=8
.ends
*
* File: G3_AND2_N2.pex.netlist
* Created: Mon Feb 28 10:46:36 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_AND2_N2_VSS 2 3 5 6 8 9 11 13 27 28 30 49 62 67 73 78 83 88 97 102
+ 111 112 116 117 122 128 130 135 136 137 139 Vss
c70 137 Vss 3.78257e-19
c71 136 Vss 3.62111e-19
c72 135 Vss 0.00438377f
c73 130 Vss 0.00256681f
c74 128 Vss 0.00549491f
c75 122 Vss 0.00414054f
c76 117 Vss 8.38241e-19
c77 116 Vss 0.00175385f
c78 112 Vss 7.28672e-19
c79 111 Vss 0.00525523f
c80 102 Vss 0.00402938f
c81 97 Vss 0.00450731f
c82 88 Vss 7.10513e-22
c83 83 Vss 4.8239e-19
c84 78 Vss 0.00106653f
c85 73 Vss 0.00125808f
c86 67 Vss 0.00537538f
c87 62 Vss 0.00490594f
c88 58 Vss 0.0299355f
c89 57 Vss 0.0299355f
c90 50 Vss 0.0347118f
c91 49 Vss 0.0994217f
c92 41 Vss 0.106723f
c93 35 Vss 0.0688517f
c94 30 Vss 5.38535e-20
c95 28 Vss 0.0340588f
c96 27 Vss 0.064644f
c97 11 Vss 0.134525f
c98 9 Vss 0.134971f
c99 8 Vss 0.133544f
c100 6 Vss 0.134177f
c101 5 Vss 0.138048f
c102 3 Vss 0.135913f
r103 135 139 0.326018
r104 134 135 5.08479
r105 130 134 0.655813
r106 129 137 0.494161
r107 128 139 0.326018
r108 128 129 10.1279
r109 124 137 0.128424
r110 123 136 0.494161
r111 122 137 0.494161
r112 122 123 10.378
r113 118 136 0.128424
r114 116 136 0.494161
r115 116 117 4.33457
r116 111 117 0.652036
r117 110 112 0.655813
r118 110 111 16.6297
r119 88 130 1.82344
r120 83 102 1.16709
r121 83 124 2.66743
r122 78 97 1.16709
r123 78 118 2.16729
r124 73 112 1.82344
r125 67 88 1.16709
r126 62 73 1.16709
r127 52 102 0.0476429
r128 50 52 1.45875
r129 49 53 0.652036
r130 49 52 1.45875
r131 46 50 0.652036
r132 42 58 0.494161
r133 41 43 0.652036
r134 41 42 2.9175
r135 37 58 0.128424
r136 36 57 0.494161
r137 35 58 0.494161
r138 35 36 2.8008
r139 31 57 0.128424
r140 30 97 0.238214
r141 28 30 1.4004
r142 27 57 0.494161
r143 27 30 1.5171
r144 24 28 0.652036
r145 13 67 0.185659
r146 11 46 3.8511
r147 9 53 3.8511
r148 8 43 3.8511
r149 6 37 3.8511
r150 5 24 3.8511
r151 3 31 3.8511
r152 2 62 0.185659
.ends

.subckt PM_G3_AND2_N2_VDD 1 3 5 7 8 10 24 26 33 43 48 53 55 56 60 62 63 66 70 72
+ 74 76 78 79 81 87 96 Vss
c85 96 Vss 0.00462548f
c86 87 Vss 0.00521601f
c87 79 Vss 4.60053e-19
c88 78 Vss 4.52364e-19
c89 76 Vss 0.00122604f
c90 74 Vss 6.12561e-19
c91 72 Vss 0.00375739f
c92 70 Vss 0.001382f
c93 66 Vss 0.00251556f
c94 63 Vss 8.66752e-19
c95 62 Vss 0.00754689f
c96 60 Vss 0.0017718f
c97 57 Vss 0.00173794f
c98 56 Vss 0.010708f
c99 55 Vss 0.00235908f
c100 53 Vss 0.00679887f
c101 48 Vss 0.00711219f
c102 43 Vss 0.00386059f
c103 33 Vss 0.0357726f
c104 32 Vss 0.102409f
c105 26 Vss 0.170515f
c106 24 Vss 0.0339269f
c107 10 Vss 0.136393f
c108 8 Vss 0.13497f
c109 7 Vss 0.00143442f
c110 1 Vss 0.117228f
r111 76 96 1.16709
r112 74 81 0.326018
r113 74 76 2.66743
r114 73 79 0.494161
r115 72 81 0.326018
r116 72 73 7.46046
r117 68 79 0.128424
r118 68 70 5.75164
r119 66 87 1.16709
r120 64 66 3.83443
r121 62 79 0.494161
r122 62 63 13.0037
r123 58 78 0.0828784
r124 58 60 1.82344
r125 56 64 0.652036
r126 56 57 10.0862
r127 55 63 0.652036
r128 54 78 0.551426
r129 54 55 5.08479
r130 53 78 0.551426
r131 52 57 0.652036
r132 52 53 13.0454
r133 48 70 1.16709
r134 43 60 1.16709
r135 35 96 0.0476429
r136 33 35 1.45875
r137 32 36 0.652036
r138 32 35 1.45875
r139 28 33 0.652036
r140 26 87 0.428786
r141 24 26 5.3682
r142 20 24 0.652036
r143 10 36 3.8511
r144 8 28 3.8511
r145 7 48 0.185659
r146 5 48 0.185659
r147 3 43 0.185659
r148 1 20 3.1509
.ends

.subckt PM_G3_AND2_N2_A 2 4 10 13 18 21 26 31 Vss
c26 31 Vss 0.00351072f
c27 26 Vss 0.00323449f
c28 18 Vss 9.2489e-19
c29 13 Vss 0.112394f
c30 2 Vss 0.112081f
r31 23 31 1.16709
r32 21 23 2.95918
r33 18 26 1.16709
r34 18 21 2.41736
r35 13 31 0.50025
r36 10 26 0.50025
r37 4 13 3.09255
r38 2 10 3.09255
.ends

.subckt PM_G3_AND2_N2_NET1 2 4 6 8 10 24 27 38 42 46 50 52 56 68 Vss
c52 68 Vss 0.00584624f
c53 58 Vss 1.47786e-19
c54 56 Vss 0.00230674f
c55 52 Vss 0.00700301f
c56 50 Vss 0.00103961f
c57 46 Vss 7.16542e-19
c58 42 Vss 0.00585482f
c59 38 Vss 0.00349773f
c60 27 Vss 9.81095e-20
c61 24 Vss 0.227317f
c62 21 Vss 0.125908f
c63 19 Vss 0.0247918f
c64 10 Vss 0.139046f
c65 6 Vss 0.00143442f
r66 56 68 1.16709
r67 54 56 3.45932
r68 53 58 0.128424
r69 52 54 0.652036
r70 52 53 7.46046
r71 48 58 0.494161
r72 48 50 6.54354
r73 44 58 0.494161
r74 44 46 3.83443
r75 42 50 1.16709
r76 38 46 1.16709
r77 27 68 0.0476429
r78 25 27 0.326018
r79 25 27 0.1167
r80 24 28 0.652036
r81 24 27 6.7686
r82 21 68 0.357321
r83 19 27 0.326018
r84 19 21 0.40845
r85 10 28 3.8511
r86 8 21 3.44265
r87 6 42 0.185659
r88 4 42 0.185659
r89 2 38 0.185659
.ends

.subckt PM_G3_AND2_N2_B 2 4 10 11 14 21 Vss
c26 21 Vss 3.50736e-19
c27 14 Vss 0.181075f
c28 11 Vss 0.0348746f
c29 10 Vss 0.288064f
c30 2 Vss 0.277377f
r31 18 21 0.0729375
r32 14 18 1.16709
r33 12 14 2.1006
r34 10 12 0.652036
r35 10 11 8.92755
r36 7 11 0.652036
r37 4 14 4.3179
r38 2 7 8.57745
.ends

.subckt PM_G3_AND2_N2_Z 2 4 13 18 Vss
c13 13 Vss 0.0052353f
c14 4 Vss 0.00143442f
r15 13 18 1.16709
r16 4 13 0.185659
r17 2 13 0.185659
.ends

.subckt G3_AND2_N2  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI5.X0 N_NET1_XI5.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_B_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW8
XI10.X0 N_NET1_XI10.X0_D N_VSS_XI10.X0_PGD N_A_XI10.X0_CG N_VSS_XI10.X0_PGS
+ N_VDD_XI10.X0_S TIGFET_HPNW8
XI6.X0 N_NET1_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGS
+ N_VDD_XI6.X0_S TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VSS_XI4.X0_PGD N_NET1_XI4.X0_CG N_VSS_XI4.X0_PGS
+ N_VDD_XI4.X0_S TIGFET_HPNW8
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_NET1_XI3.X0_CG N_VDD_XI3.X0_PGS
+ N_VSS_XI3.X0_S TIGFET_HPNW8
*
x_PM_G3_AND2_N2_VSS N_VSS_XI5.X0_S N_VSS_XI10.X0_PGD N_VSS_XI10.X0_PGS
+ N_VSS_XI6.X0_PGD N_VSS_XI6.X0_PGS N_VSS_XI4.X0_PGD N_VSS_XI4.X0_PGS
+ N_VSS_XI3.X0_S N_VSS_c_13_p N_VSS_c_14_p N_VSS_c_46_p N_VSS_c_2_p N_VSS_c_3_p
+ N_VSS_c_65_p N_VSS_c_4_p N_VSS_c_8_p N_VSS_c_24_p N_VSS_c_66_p N_VSS_c_9_p
+ N_VSS_c_26_p N_VSS_c_5_p N_VSS_c_6_p N_VSS_c_17_p N_VSS_c_20_p N_VSS_c_18_p
+ N_VSS_c_32_p N_VSS_c_70_p N_VSS_c_37_p N_VSS_c_19_p N_VSS_c_33_p VSS Vss
+ PM_G3_AND2_N2_VSS
x_PM_G3_AND2_N2_VDD N_VDD_XI5.X0_PGD N_VDD_XI10.X0_S N_VDD_XI6.X0_S
+ N_VDD_XI4.X0_S N_VDD_XI3.X0_PGD N_VDD_XI3.X0_PGS N_VDD_c_148_p N_VDD_c_130_p
+ N_VDD_c_72_n N_VDD_c_125_p N_VDD_c_126_p N_VDD_c_73_n N_VDD_c_77_n
+ N_VDD_c_81_n N_VDD_c_82_n N_VDD_c_83_n N_VDD_c_90_n N_VDD_c_123_p N_VDD_c_91_n
+ N_VDD_c_98_n N_VDD_c_104_n N_VDD_c_105_n N_VDD_c_108_n N_VDD_c_109_n VDD
+ N_VDD_c_119_p N_VDD_c_110_n Vss PM_G3_AND2_N2_VDD
x_PM_G3_AND2_N2_A N_A_XI5.X0_CG N_A_XI10.X0_CG N_A_c_164_n N_A_c_156_n
+ N_A_c_157_n A N_A_c_167_n N_A_c_160_n Vss PM_G3_AND2_N2_A
x_PM_G3_AND2_N2_NET1 N_NET1_XI5.X0_D N_NET1_XI10.X0_D N_NET1_XI6.X0_D
+ N_NET1_XI4.X0_CG N_NET1_XI3.X0_CG N_NET1_c_182_n N_NET1_c_183_n N_NET1_c_184_n
+ N_NET1_c_199_n N_NET1_c_186_n N_NET1_c_189_n N_NET1_c_190_n N_NET1_c_191_n
+ N_NET1_c_193_n Vss PM_G3_AND2_N2_NET1
x_PM_G3_AND2_N2_B N_B_XI5.X0_PGS N_B_XI6.X0_CG N_B_c_234_n N_B_c_236_n
+ N_B_c_241_n B Vss PM_G3_AND2_N2_B
x_PM_G3_AND2_N2_Z N_Z_XI4.X0_D N_Z_XI3.X0_D N_Z_c_260_n Z Vss PM_G3_AND2_N2_Z
cc_1 N_VSS_XI4.X0_PGD N_VDD_XI3.X0_PGD 0.00195824f
cc_2 N_VSS_c_2_p N_VDD_c_72_n 0.00195824f
cc_3 N_VSS_c_3_p N_VDD_c_73_n 9.5668e-19
cc_4 N_VSS_c_4_p N_VDD_c_73_n 0.00165395f
cc_5 N_VSS_c_5_p N_VDD_c_73_n 0.00670587f
cc_6 N_VSS_c_6_p N_VDD_c_73_n 0.00189531f
cc_7 N_VSS_XI10.X0_PGS N_VDD_c_77_n 2.75457e-19
cc_8 N_VSS_c_8_p N_VDD_c_77_n 4.50283e-19
cc_9 N_VSS_c_9_p N_VDD_c_77_n 3.70842e-19
cc_10 N_VSS_c_5_p N_VDD_c_77_n 0.00345577f
cc_11 N_VSS_c_4_p N_VDD_c_81_n 0.00247496f
cc_12 N_VSS_c_4_p N_VDD_c_82_n 4.32396e-19
cc_13 N_VSS_c_13_p N_VDD_c_83_n 0.00151774f
cc_14 N_VSS_c_14_p N_VDD_c_83_n 3.51214e-19
cc_15 N_VSS_c_8_p N_VDD_c_83_n 0.00161703f
cc_16 N_VSS_c_9_p N_VDD_c_83_n 2.03837e-19
cc_17 N_VSS_c_17_p N_VDD_c_83_n 0.00348097f
cc_18 N_VSS_c_18_p N_VDD_c_83_n 0.0059139f
cc_19 N_VSS_c_19_p N_VDD_c_83_n 7.61747e-19
cc_20 N_VSS_c_20_p N_VDD_c_90_n 0.00107346f
cc_21 N_VSS_XI6.X0_PGS N_VDD_c_91_n 2.23834e-19
cc_22 N_VSS_XI4.X0_PGS N_VDD_c_91_n 2.29703e-19
cc_23 N_VSS_c_8_p N_VDD_c_91_n 6.50938e-19
cc_24 N_VSS_c_24_p N_VDD_c_91_n 0.00193467f
cc_25 N_VSS_c_9_p N_VDD_c_91_n 2.56577e-19
cc_26 N_VSS_c_26_p N_VDD_c_91_n 9.55109e-19
cc_27 N_VSS_c_5_p N_VDD_c_91_n 3.54686e-19
cc_28 N_VSS_c_2_p N_VDD_c_98_n 4.82224e-19
cc_29 N_VSS_c_24_p N_VDD_c_98_n 0.00118142f
cc_30 N_VSS_c_26_p N_VDD_c_98_n 2.13453e-19
cc_31 N_VSS_c_18_p N_VDD_c_98_n 0.00133442f
cc_32 N_VSS_c_32_p N_VDD_c_98_n 0.00433318f
cc_33 N_VSS_c_33_p N_VDD_c_98_n 8.13487e-19
cc_34 N_VSS_c_32_p N_VDD_c_104_n 0.00157826f
cc_35 N_VSS_c_24_p N_VDD_c_105_n 9.21598e-19
cc_36 N_VSS_c_26_p N_VDD_c_105_n 3.82294e-19
cc_37 N_VSS_c_37_p N_VDD_c_105_n 5.22507e-19
cc_38 N_VSS_c_5_p N_VDD_c_108_n 0.00100712f
cc_39 N_VSS_c_18_p N_VDD_c_109_n 9.86755e-19
cc_40 N_VSS_c_24_p N_VDD_c_110_n 3.48267e-19
cc_41 N_VSS_c_26_p N_VDD_c_110_n 6.46219e-19
cc_42 N_VSS_c_9_p N_A_c_156_n 0.00249847f
cc_43 N_VSS_c_8_p N_A_c_157_n 2.94885e-19
cc_44 N_VSS_c_9_p N_A_c_157_n 3.71222e-19
cc_45 N_VSS_c_5_p N_A_c_157_n 0.00147463f
cc_46 N_VSS_c_46_p N_A_c_160_n 3.96531e-19
cc_47 N_VSS_c_8_p N_A_c_160_n 2.87758e-19
cc_48 N_VSS_c_9_p N_A_c_160_n 8.98435e-19
cc_49 N_VSS_XI4.X0_PGD N_NET1_c_182_n 4.26252e-19
cc_50 N_VSS_c_26_p N_NET1_c_183_n 9.4551e-19
cc_51 N_VSS_c_3_p N_NET1_c_184_n 3.43419e-19
cc_52 N_VSS_c_4_p N_NET1_c_184_n 3.48267e-19
cc_53 N_VSS_c_3_p N_NET1_c_186_n 3.48267e-19
cc_54 N_VSS_c_4_p N_NET1_c_186_n 8.50248e-19
cc_55 N_VSS_c_5_p N_NET1_c_186_n 5.59972e-19
cc_56 N_VSS_c_18_p N_NET1_c_189_n 2.3523e-19
cc_57 N_VSS_c_18_p N_NET1_c_190_n 4.47676e-19
cc_58 N_VSS_c_24_p N_NET1_c_191_n 5.58211e-19
cc_59 N_VSS_c_26_p N_NET1_c_191_n 3.49408e-19
cc_60 N_VSS_c_24_p N_NET1_c_193_n 3.2351e-19
cc_61 N_VSS_c_26_p N_NET1_c_193_n 2.68747e-19
cc_62 N_VSS_XI10.X0_PGD N_B_c_234_n 8.28117e-19
cc_63 N_VSS_XI6.X0_PGD N_B_c_234_n 8.28117e-19
cc_64 N_VSS_XI10.X0_PGS N_B_c_236_n 9.94582e-19
cc_65 N_VSS_c_65_p N_Z_c_260_n 3.43419e-19
cc_66 N_VSS_c_66_p N_Z_c_260_n 3.48267e-19
cc_67 N_VSS_c_65_p Z 3.48267e-19
cc_68 N_VSS_c_66_p Z 4.99861e-19
cc_69 N_VSS_c_32_p Z 2.34298e-19
cc_70 N_VSS_c_70_p Z 2.7826e-19
cc_71 N_VDD_XI5.X0_PGD N_A_XI5.X0_CG 5.26351e-19
cc_72 N_VDD_c_81_n N_A_c_164_n 3.14632e-19
cc_73 N_VDD_c_73_n N_A_c_157_n 0.00285022f
cc_74 N_VDD_c_81_n N_A_c_157_n 5.83159e-19
cc_75 N_VDD_XI5.X0_PGD N_A_c_167_n 2.78309e-19
cc_76 N_VDD_c_73_n N_A_c_167_n 3.66936e-19
cc_77 N_VDD_c_81_n N_A_c_167_n 3.4118e-19
cc_78 N_VDD_c_119_p N_A_c_167_n 4.44265e-19
cc_79 N_VDD_c_73_n N_A_c_160_n 4.70132e-19
cc_80 N_VDD_XI3.X0_PGD N_NET1_c_182_n 4.29017e-19
cc_81 N_VDD_c_81_n N_NET1_c_184_n 9.18655e-19
cc_82 N_VDD_c_123_p N_NET1_c_184_n 8.835e-19
cc_83 N_VDD_c_119_p N_NET1_c_184_n 0.00132057f
cc_84 N_VDD_c_125_p N_NET1_c_199_n 3.43419e-19
cc_85 N_VDD_c_126_p N_NET1_c_199_n 3.43419e-19
cc_86 N_VDD_c_82_n N_NET1_c_199_n 3.72199e-19
cc_87 N_VDD_c_83_n N_NET1_c_199_n 3.02646e-19
cc_88 N_VDD_c_91_n N_NET1_c_199_n 3.48267e-19
cc_89 N_VDD_c_130_p N_NET1_c_186_n 7.85476e-19
cc_90 N_VDD_c_73_n N_NET1_c_186_n 9.00704e-19
cc_91 N_VDD_c_81_n N_NET1_c_186_n 0.00168791f
cc_92 N_VDD_c_123_p N_NET1_c_186_n 0.00355804f
cc_93 N_VDD_c_119_p N_NET1_c_186_n 8.835e-19
cc_94 N_VDD_c_125_p N_NET1_c_189_n 3.48267e-19
cc_95 N_VDD_c_126_p N_NET1_c_189_n 3.48267e-19
cc_96 N_VDD_c_82_n N_NET1_c_189_n 8.08807e-19
cc_97 N_VDD_c_83_n N_NET1_c_189_n 4.24175e-19
cc_98 N_VDD_c_91_n N_NET1_c_189_n 7.1497e-19
cc_99 N_VDD_c_130_p N_NET1_c_190_n 3.97408e-19
cc_100 N_VDD_c_126_p N_NET1_c_190_n 2.52932e-19
cc_101 N_VDD_c_123_p N_NET1_c_190_n 0.001476f
cc_102 N_VDD_c_91_n N_NET1_c_190_n 5.44012e-19
cc_103 N_VDD_c_119_p N_NET1_c_190_n 0.00114101f
cc_104 N_VDD_XI5.X0_PGD N_B_XI5.X0_PGS 0.00153355f
cc_105 N_VDD_c_73_n N_B_XI5.X0_PGS 7.45044e-19
cc_106 N_VDD_c_81_n N_B_XI5.X0_PGS 3.02077e-19
cc_107 N_VDD_c_148_p N_B_c_234_n 0.00419437f
cc_108 N_VDD_c_119_p N_B_c_241_n 7.17663e-19
cc_109 N_VDD_c_126_p N_Z_c_260_n 3.43419e-19
cc_110 N_VDD_c_91_n N_Z_c_260_n 3.48267e-19
cc_111 N_VDD_c_98_n N_Z_c_260_n 3.02646e-19
cc_112 N_VDD_c_126_p Z 3.48267e-19
cc_113 N_VDD_c_91_n Z 7.09569e-19
cc_114 N_VDD_c_98_n Z 4.04319e-19
cc_115 N_A_c_157_n N_NET1_c_186_n 0.00799902f
cc_116 N_A_c_167_n N_NET1_c_186_n 8.66889e-19
cc_117 N_A_c_160_n N_NET1_c_189_n 9.68342e-19
cc_118 N_A_XI5.X0_CG N_B_XI5.X0_PGS 4.87172e-19
cc_119 N_A_c_157_n N_B_XI5.X0_PGS 4.74011e-19
cc_120 N_A_c_167_n N_B_XI5.X0_PGS 5.6636e-19
cc_121 N_A_c_157_n N_B_c_234_n 2.0632e-19
cc_122 N_A_c_167_n N_B_c_234_n 7.2846e-19
cc_123 N_A_c_160_n N_B_c_234_n 0.00228839f
cc_124 N_A_c_160_n N_B_c_241_n 9.27569e-19
cc_125 N_NET1_c_199_n N_B_c_234_n 3.74089e-19
cc_126 N_NET1_c_189_n N_B_c_234_n 3.943e-19
cc_127 N_NET1_c_190_n N_B_c_234_n 2.82146e-19
cc_128 N_NET1_c_189_n N_B_c_241_n 0.00116203f
cc_129 N_NET1_c_190_n N_B_c_241_n 5.60175e-19
cc_130 N_NET1_c_191_n N_B_c_241_n 3.86148e-19
cc_131 N_NET1_c_193_n N_B_c_241_n 0.00196155f
cc_132 N_NET1_c_189_n B 0.00147455f
cc_133 N_NET1_c_190_n B 8.26881e-19
cc_134 N_NET1_c_191_n B 5.75904e-19
cc_135 N_NET1_c_193_n B 3.48267e-19
cc_136 N_NET1_c_182_n N_Z_c_260_n 6.55689e-19
*
.ends
*
*
.subckt AND2_HPNW8 A B Y VDD VSS
xgate (VSS VDD A B Y) G3_AND2_N2
.ends
*
* File: G2_AOI21_N2.pex.netlist
* Created: Mon Apr 11 18:40:10 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_AOI21_N2_VSS 2 4 6 8 19 30 35 38 43 48 57 66 67 69 77 78 79 84 86
+ 88 89 Vss
c51 89 Vss 4.28045e-19
c52 86 Vss 0.00486026f
c53 84 Vss 0.00155386f
c54 79 Vss 0.00128356f
c55 78 Vss 4.65637e-19
c56 77 Vss 0.00250049f
c57 69 Vss 0.00102564f
c58 67 Vss 0.00986383f
c59 66 Vss 0.00273179f
c60 65 Vss 0.00133186f
c61 57 Vss 0.00579208f
c62 48 Vss 2.73256e-19
c63 43 Vss 0.00178422f
c64 38 Vss 0.00142279f
c65 35 Vss 0.00389683f
c66 30 Vss 0.00549227f
c67 25 Vss 0.0828998f
c68 19 Vss 0.0350566f
c69 18 Vss 0.0688416f
c70 8 Vss 0.135691f
c71 4 Vss 0.134006f
r72 85 89 0.551426
r73 85 86 15.5878
r74 84 89 0.551426
r75 83 84 4.58464
r76 79 89 0.0828784
r77 77 86 0.652036
r78 77 78 4.33457
r79 73 78 0.652036
r80 68 88 0.326018
r81 67 83 0.652036
r82 67 68 15.6711
r83 66 69 0.655813
r84 65 88 0.326018
r85 65 66 4.58464
r86 48 79 1.82344
r87 43 57 1.16709
r88 43 73 2.16729
r89 38 69 1.82344
r90 35 48 1.16709
r91 30 38 1.16709
r92 25 57 0.0476429
r93 23 25 2.04225
r94 20 23 0.0685365
r95 18 23 0.5835
r96 18 19 2.8008
r97 15 19 0.652036
r98 8 20 3.8511
r99 6 35 0.185659
r100 4 15 3.8511
r101 2 30 0.185659
.ends

.subckt PM_G2_AOI21_N2_VDD 2 4 6 8 10 29 37 42 45 46 48 50 54 56 57 58 62 63 65
+ 67 68 74 Vss
c58 74 Vss 0.00462133f
c59 68 Vss 4.52364e-19
c60 65 Vss 0.00203839f
c61 63 Vss 0.00821501f
c62 62 Vss 8.61193e-19
c63 58 Vss 0.00179763f
c64 57 Vss 6.04409e-19
c65 56 Vss 0.00220637f
c66 54 Vss 0.00139836f
c67 51 Vss 0.00169975f
c68 50 Vss 0.0126653f
c69 48 Vss 0.00162243f
c70 46 Vss 0.00140335f
c71 45 Vss 0.00324454f
c72 42 Vss 0.00402078f
c73 37 Vss 0.00544429f
c74 33 Vss 0.0307649f
c75 29 Vss 1.05042e-19
c76 26 Vss 0.101606f
c77 22 Vss 0.035898f
c78 21 Vss 0.0712517f
c79 8 Vss 0.135377f
c80 6 Vss 0.136126f
c81 2 Vss 0.135008f
r82 64 68 0.551426
r83 64 65 4.58464
r84 63 68 0.551426
r85 62 67 0.326018
r86 62 63 15.5878
r87 58 68 0.0828784
r88 58 60 1.82344
r89 56 67 0.326018
r90 56 57 4.37625
r91 54 74 1.16709
r92 52 57 0.652036
r93 52 54 2.16729
r94 50 65 0.652036
r95 50 51 15.7128
r96 46 48 1.85991
r97 45 51 0.652036
r98 44 46 0.655813
r99 44 45 4.58464
r100 42 60 1.16709
r101 37 48 1.16709
r102 29 74 0.0476429
r103 27 33 0.494161
r104 27 29 1.45875
r105 26 30 0.652036
r106 26 29 1.45875
r107 23 33 0.128424
r108 21 33 0.494161
r109 21 22 2.8008
r110 18 22 0.652036
r111 10 42 0.185659
r112 8 30 3.8511
r113 6 23 3.8511
r114 4 37 0.185659
r115 2 18 3.8511
.ends

.subckt PM_G2_AOI21_N2_B 2 4 20 25 28 Vss
c17 28 Vss 0.00498247f
c18 25 Vss 6.10536e-19
c19 20 Vss 0.0915067f
c20 16 Vss 0.0598477f
c21 4 Vss 0.157143f
c22 2 Vss 0.372582f
r23 25 28 1.16709
r24 18 20 2.04225
r25 16 28 0.197068
r26 13 16 1.2837
r27 10 20 0.0685365
r28 8 18 0.0685365
r29 7 13 0.0685365
r30 4 10 4.3179
r31 2 8 9.9195
r32 2 7 3.8511
.ends

.subckt PM_G2_AOI21_N2_C 2 4 6 17 24 28 31 34 38 43 56 Vss
c46 56 Vss 0.00123749f
c47 43 Vss 0.0052622f
c48 38 Vss 0.00284502f
c49 34 Vss 0.00609886f
c50 28 Vss 0.0947914f
c51 24 Vss 0.0843207f
c52 17 Vss 3.53906e-19
c53 6 Vss 0.232307f
c54 4 Vss 0.201668f
c55 2 Vss 0.134559f
r56 52 56 0.652036
r57 38 56 5.16814
r58 34 43 1.16709
r59 34 52 10.4196
r60 31 34 0.145875
r61 26 28 2.04225
r62 24 43 0.0476429
r63 21 24 1.92555
r64 18 28 0.0685365
r65 17 38 1.16709
r66 13 26 0.0685365
r67 13 17 2.8008
r68 10 21 0.0685365
r69 6 18 7.1187
r70 4 17 4.3179
r71 2 10 3.8511
.ends

.subckt PM_G2_AOI21_N2_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00256251f
c33 27 Vss 0.00470045f
c34 23 Vss 0.00695334f
c35 8 Vss 0.00143442f
c36 6 Vss 0.00143442f
r37 33 35 7.002
r38 30 33 4.00114
r39 27 35 1.16709
r40 23 30 1.16709
r41 8 27 0.185659
r42 6 23 0.185659
r43 4 27 0.185659
r44 2 23 0.185659
.ends

.subckt PM_G2_AOI21_N2_A 2 4 10 11 13 14 15 20 24 29 32 Vss
c34 32 Vss 9.11501e-19
c35 29 Vss 4.23286e-19
c36 24 Vss 1.80739e-19
c37 20 Vss 0.136821f
c38 18 Vss 0.0247918f
c39 15 Vss 0.0322409f
c40 14 Vss 0.0730777f
c41 13 Vss 0.0312529f
c42 11 Vss 0.0324953f
c43 10 Vss 0.122088f
c44 2 Vss 0.238343f
r45 26 32 1.16709
r46 26 29 0.0729375
r47 24 32 0.262036
r48 20 32 0.238214
r49 18 24 0.326018
r50 18 20 0.64185
r51 15 24 2.50905
r52 14 24 0.326018
r53 14 24 0.1167
r54 13 15 0.652036
r55 12 13 1.22535
r56 10 12 0.652036
r57 10 11 3.09255
r58 7 11 0.652036
r59 4 20 3.7344
r60 2 7 7.4688
.ends

.subckt G2_AOI21_N2  VSS VDD B C Z A
*
* A	A
* Z	Z
* C	C
* B	B
* VDD	VDD
* VSS	VSS
XI14.X0 N_Z_XI14.X0_D N_VDD_XI14.X0_PGD N_A_XI14.X0_CG N_B_XI14.X0_PGS
+ N_VSS_XI14.X0_S TIGFET_HPNW8
XI12.X0 N_Z_XI12.X0_D N_VSS_XI12.X0_PGD N_B_XI12.X0_CG N_C_XI12.X0_PGS
+ N_VDD_XI12.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_VDD_XI15.X0_PGD N_C_XI15.X0_CG N_VDD_XI15.X0_PGS
+ N_VSS_XI15.X0_S TIGFET_HPNW8
XI13.X0 N_Z_XI13.X0_D N_VSS_XI13.X0_PGD N_A_XI13.X0_CG N_C_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW8
*
x_PM_G2_AOI21_N2_VSS N_VSS_XI14.X0_S N_VSS_XI12.X0_PGD N_VSS_XI15.X0_S
+ N_VSS_XI13.X0_PGD N_VSS_c_3_p N_VSS_c_35_p N_VSS_c_8_p N_VSS_c_2_p N_VSS_c_4_p
+ N_VSS_c_9_p N_VSS_c_5_p N_VSS_c_22_p N_VSS_c_10_p N_VSS_c_1_p N_VSS_c_6_p
+ N_VSS_c_7_p N_VSS_c_12_p N_VSS_c_15_p N_VSS_c_16_p VSS N_VSS_c_17_p Vss
+ PM_G2_AOI21_N2_VSS
x_PM_G2_AOI21_N2_VDD N_VDD_XI14.X0_PGD N_VDD_XI12.X0_S N_VDD_XI15.X0_PGD
+ N_VDD_XI15.X0_PGS N_VDD_XI13.X0_S N_VDD_c_80_p N_VDD_c_95_p N_VDD_c_96_p
+ N_VDD_c_79_p N_VDD_c_52_n N_VDD_c_53_n N_VDD_c_54_n N_VDD_c_74_p N_VDD_c_59_n
+ N_VDD_c_62_n N_VDD_c_63_n N_VDD_c_64_n N_VDD_c_65_n N_VDD_c_69_n VDD
+ N_VDD_c_72_n N_VDD_c_75_p Vss PM_G2_AOI21_N2_VDD
x_PM_G2_AOI21_N2_B N_B_XI14.X0_PGS N_B_XI12.X0_CG N_B_c_118_p B N_B_c_115_n Vss
+ PM_G2_AOI21_N2_B
x_PM_G2_AOI21_N2_C N_C_XI12.X0_PGS N_C_XI15.X0_CG N_C_XI13.X0_PGS N_C_c_139_n
+ N_C_c_142_n N_C_c_143_n C N_C_c_128_n N_C_c_131_n N_C_c_132_n N_C_c_136_n Vss
+ PM_G2_AOI21_N2_C
x_PM_G2_AOI21_N2_Z N_Z_XI14.X0_D N_Z_XI12.X0_D N_Z_XI15.X0_D N_Z_XI13.X0_D
+ N_Z_c_173_n N_Z_c_183_n N_Z_c_177_n Z Vss PM_G2_AOI21_N2_Z
x_PM_G2_AOI21_N2_A N_A_XI14.X0_CG N_A_XI13.X0_CG N_A_c_205_n N_A_c_217_n
+ N_A_c_218_n N_A_c_206_n N_A_c_219_n N_A_c_225_n N_A_c_207_n A N_A_c_210_n Vss
+ PM_G2_AOI21_N2_A
cc_1 N_VSS_c_1_p N_VDD_c_52_n 3.73937e-19
cc_2 N_VSS_c_2_p N_VDD_c_53_n 5.43852e-19
cc_3 N_VSS_c_3_p N_VDD_c_54_n 0.0012732f
cc_4 N_VSS_c_4_p N_VDD_c_54_n 0.00161703f
cc_5 N_VSS_c_5_p N_VDD_c_54_n 2.26455e-19
cc_6 N_VSS_c_6_p N_VDD_c_54_n 0.00447304f
cc_7 N_VSS_c_7_p N_VDD_c_54_n 0.00169823f
cc_8 N_VSS_c_8_p N_VDD_c_59_n 3.4118e-19
cc_9 N_VSS_c_9_p N_VDD_c_59_n 4.19648e-19
cc_10 N_VSS_c_10_p N_VDD_c_59_n 0.00353938f
cc_11 N_VSS_c_10_p N_VDD_c_62_n 0.00161744f
cc_12 N_VSS_c_12_p N_VDD_c_63_n 4.54377e-19
cc_13 N_VSS_c_10_p N_VDD_c_64_n 0.00106833f
cc_14 N_VSS_c_9_p N_VDD_c_65_n 0.00187494f
cc_15 N_VSS_c_15_p N_VDD_c_65_n 0.00340036f
cc_16 N_VSS_c_16_p N_VDD_c_65_n 0.00745699f
cc_17 N_VSS_c_17_p N_VDD_c_65_n 9.16632e-19
cc_18 N_VSS_c_4_p N_VDD_c_69_n 4.42007e-19
cc_19 N_VSS_c_5_p N_VDD_c_69_n 4.06699e-19
cc_20 N_VSS_c_16_p N_VDD_c_69_n 0.00303867f
cc_21 N_VSS_c_16_p N_VDD_c_72_n 0.00115015f
cc_22 N_VSS_c_22_p B 3.69138e-19
cc_23 N_VSS_c_10_p B 3.52052e-19
cc_24 N_VSS_XI12.X0_PGD N_C_XI12.X0_PGS 0.00151939f
cc_25 N_VSS_c_4_p N_C_c_128_n 8.90801e-19
cc_26 N_VSS_c_5_p N_C_c_128_n 3.44698e-19
cc_27 N_VSS_c_16_p N_C_c_128_n 0.00169235f
cc_28 N_VSS_c_16_p N_C_c_131_n 5.11302e-19
cc_29 N_VSS_XI12.X0_PGD N_C_c_132_n 3.23173e-19
cc_30 N_VSS_c_3_p N_C_c_132_n 0.00480946f
cc_31 N_VSS_c_4_p N_C_c_132_n 3.44698e-19
cc_32 N_VSS_c_5_p N_C_c_132_n 6.61756e-19
cc_33 N_VSS_c_10_p N_C_c_136_n 0.00251881f
cc_34 N_VSS_c_16_p N_C_c_136_n 3.90377e-19
cc_35 N_VSS_c_35_p N_Z_c_173_n 3.43419e-19
cc_36 N_VSS_c_8_p N_Z_c_173_n 3.43419e-19
cc_37 N_VSS_c_2_p N_Z_c_173_n 3.48267e-19
cc_38 N_VSS_c_9_p N_Z_c_173_n 3.48267e-19
cc_39 N_VSS_c_35_p N_Z_c_177_n 3.48267e-19
cc_40 N_VSS_c_8_p N_Z_c_177_n 3.48267e-19
cc_41 N_VSS_c_2_p N_Z_c_177_n 5.71987e-19
cc_42 N_VSS_c_9_p N_Z_c_177_n 5.71987e-19
cc_43 N_VSS_c_10_p N_Z_c_177_n 3.08274e-19
cc_44 N_VSS_c_16_p N_Z_c_177_n 7.49935e-19
cc_45 N_VSS_XI12.X0_PGD N_A_c_205_n 7.49544e-19
cc_46 N_VSS_XI13.X0_PGD N_A_c_206_n 0.00161855f
cc_47 N_VSS_c_5_p N_A_c_207_n 9.11194e-19
cc_48 N_VSS_c_4_p A 3.22909e-19
cc_49 N_VSS_c_5_p A 3.2351e-19
cc_50 N_VSS_c_4_p N_A_c_210_n 3.2351e-19
cc_51 N_VSS_c_5_p N_A_c_210_n 2.68747e-19
cc_52 N_VDD_XI14.X0_PGD N_B_XI14.X0_PGS 0.00174385f
cc_53 N_VDD_c_74_p B 6.29947e-19
cc_54 N_VDD_c_75_p B 3.48267e-19
cc_55 N_VDD_XI14.X0_PGD N_B_c_115_n 3.23173e-19
cc_56 N_VDD_c_74_p N_B_c_115_n 4.44903e-19
cc_57 N_VDD_c_75_p N_B_c_115_n 6.39485e-19
cc_58 N_VDD_c_79_p N_C_XI12.X0_PGS 2.86849e-19
cc_59 N_VDD_c_80_p N_C_c_139_n 9.37804e-19
cc_60 N_VDD_c_65_n N_C_c_139_n 5.88901e-19
cc_61 N_VDD_c_75_p N_C_c_139_n 2.68747e-19
cc_62 N_VDD_c_54_n N_C_c_142_n 3.8224e-19
cc_63 N_VDD_XI15.X0_PGS N_C_c_143_n 8.15793e-19
cc_64 N_VDD_c_65_n N_C_c_143_n 5.55843e-19
cc_65 N_VDD_c_79_p N_C_c_128_n 9.5543e-19
cc_66 N_VDD_c_53_n N_C_c_128_n 4.34676e-19
cc_67 N_VDD_c_54_n N_C_c_128_n 0.00198126f
cc_68 N_VDD_c_54_n N_C_c_131_n 6.31729e-19
cc_69 N_VDD_c_74_p N_C_c_131_n 4.21038e-19
cc_70 N_VDD_c_65_n N_C_c_131_n 4.49702e-19
cc_71 N_VDD_c_75_p N_C_c_131_n 3.2351e-19
cc_72 N_VDD_c_79_p N_C_c_132_n 3.63088e-19
cc_73 N_VDD_c_54_n N_C_c_132_n 2.64932e-19
cc_74 N_VDD_c_95_p N_Z_c_183_n 3.43419e-19
cc_75 N_VDD_c_96_p N_Z_c_183_n 3.43419e-19
cc_76 N_VDD_c_53_n N_Z_c_183_n 3.72424e-19
cc_77 N_VDD_c_54_n N_Z_c_183_n 3.4118e-19
cc_78 N_VDD_c_63_n N_Z_c_183_n 3.72199e-19
cc_79 N_VDD_c_95_p N_Z_c_177_n 3.48267e-19
cc_80 N_VDD_c_96_p N_Z_c_177_n 3.48267e-19
cc_81 N_VDD_c_53_n N_Z_c_177_n 5.09689e-19
cc_82 N_VDD_c_54_n N_Z_c_177_n 6.43655e-19
cc_83 N_VDD_c_63_n N_Z_c_177_n 7.72285e-19
cc_84 N_VDD_c_65_n N_Z_c_177_n 0.00139834f
cc_85 N_VDD_XI14.X0_PGD N_A_c_205_n 6.23873e-19
cc_86 N_VDD_XI15.X0_PGD N_A_c_206_n 3.69557e-19
cc_87 N_VDD_c_65_n A 4.8807e-19
cc_88 N_VDD_c_65_n N_A_c_210_n 3.66936e-19
cc_89 N_B_c_118_p N_C_XI12.X0_PGS 0.00196296f
cc_90 N_B_XI14.X0_PGS N_C_XI15.X0_CG 2.46172e-19
cc_91 N_B_c_118_p N_C_XI13.X0_PGS 4.66827e-19
cc_92 N_B_XI14.X0_PGS N_Z_c_177_n 2.61881e-19
cc_93 N_B_XI14.X0_PGS N_A_XI14.X0_CG 0.00881601f
cc_94 N_B_c_118_p N_A_c_217_n 0.00188162f
cc_95 N_B_XI14.X0_PGS N_A_c_218_n 6.07734e-19
cc_96 N_B_c_118_p N_A_c_219_n 0.00136534f
cc_97 N_B_c_118_p N_A_c_210_n 2.87722e-19
cc_98 N_C_c_139_n N_Z_c_177_n 9.83688e-19
cc_99 N_C_c_128_n N_Z_c_177_n 0.00274829f
cc_100 N_C_c_131_n N_Z_c_177_n 0.00329442f
cc_101 N_C_c_136_n N_Z_c_177_n 2.70867e-19
cc_102 N_C_XI15.X0_CG N_A_XI14.X0_CG 5.48933e-19
cc_103 N_C_c_139_n N_A_XI14.X0_CG 5.60239e-19
cc_104 N_C_XI13.X0_PGS N_A_c_205_n 8.10159e-19
cc_105 N_C_c_143_n N_A_c_205_n 0.00121323f
cc_106 N_C_XI13.X0_PGS N_A_c_225_n 4.5346e-19
cc_107 N_C_c_139_n N_A_c_207_n 9.47282e-19
cc_108 N_C_c_139_n A 4.56568e-19
cc_109 N_C_c_131_n A 6.34188e-19
cc_110 N_C_XI13.X0_PGS N_A_c_210_n 0.00570455f
cc_111 N_C_c_139_n N_A_c_210_n 6.1245e-19
cc_112 N_C_c_143_n N_A_c_210_n 0.00148932f
cc_113 N_C_c_131_n N_A_c_210_n 4.56568e-19
cc_114 N_Z_c_177_n N_A_XI14.X0_CG 5.52516e-19
cc_115 N_Z_c_173_n N_A_c_205_n 3.52706e-19
cc_116 N_Z_c_177_n N_A_c_205_n 3.09083e-19
cc_117 N_Z_c_183_n N_A_c_219_n 5.59623e-19
cc_118 N_Z_c_177_n A 0.00149422f
cc_119 N_Z_c_177_n N_A_c_210_n 9.63126e-19
*
.ends
*
*
.subckt AOI21_HPNW8 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 B0 Y A0) G2_AOI21_N2
.ends
*
* File: G2_BUF1_N2.pex.netlist
* Created: Wed Mar  2 15:38:39 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_BUF1_N2_VDD 2 4 7 11 28 30 32 44 48 52 54 56 57 61 65 67 71 75 78
+ 90 95 Vss
c59 95 Vss 0.0047576f
c60 90 Vss 0.00460635f
c61 80 Vss 9.22237e-19
c62 79 Vss 9.22237e-19
c63 75 Vss 0.00103298f
c64 71 Vss 9.84953e-19
c65 68 Vss 0.001766f
c66 67 Vss 0.0073616f
c67 65 Vss 0.00118372f
c68 61 Vss 0.00118372f
c69 57 Vss 0.00729501f
c70 56 Vss 0.0034296f
c71 54 Vss 0.00566164f
c72 52 Vss 0.0034296f
c73 51 Vss 0.001766f
c74 48 Vss 0.00382489f
c75 44 Vss 0.00532438f
c76 32 Vss 0.035607f
c77 31 Vss 0.102409f
c78 28 Vss 0.035607f
c79 27 Vss 0.102409f
c80 11 Vss 0.270897f
c81 7 Vss 0.270897f
r82 75 95 1.16709
r83 73 75 2.16729
r84 71 90 1.16709
r85 69 71 2.16729
r86 67 73 0.652036
r87 67 68 10.1279
r88 63 80 0.0828784
r89 63 65 1.82344
r90 59 79 0.0828784
r91 59 61 1.82344
r92 58 78 0.326018
r93 57 69 0.652036
r94 57 58 10.1279
r95 56 68 0.652036
r96 55 80 0.551426
r97 55 56 4.58464
r98 54 80 0.551426
r99 53 79 0.551426
r100 53 54 6.75193
r101 52 79 0.551426
r102 51 78 0.326018
r103 51 52 4.58464
r104 48 65 1.16709
r105 44 61 1.16709
r106 34 95 0.0476429
r107 32 34 1.45875
r108 31 38 0.652036
r109 31 34 1.45875
r110 30 90 0.0476429
r111 28 30 1.45875
r112 27 35 0.652036
r113 27 30 1.45875
r114 24 32 0.652036
r115 21 28 0.652036
r116 11 38 3.8511
r117 11 24 3.8511
r118 7 35 3.8511
r119 7 21 3.8511
r120 4 48 0.185659
r121 2 44 0.185659
.ends

.subckt PM_G2_BUF1_N2_VSS 3 7 10 12 27 28 30 31 32 45 49 52 57 62 67 72 77 97 98
+ 99 100 101 105 110 112 114 118 Vss
c56 116 Vss 6.78504e-19
c57 115 Vss 6.78504e-19
c58 114 Vss 0.00409661f
c59 112 Vss 0.00423582f
c60 110 Vss 0.0027381f
c61 105 Vss 0.0010217f
c62 101 Vss 8.62361e-19
c63 100 Vss 5.83649e-19
c64 99 Vss 0.00516968f
c65 98 Vss 5.83649e-19
c66 97 Vss 0.00631668f
c67 77 Vss 0.00400078f
c68 72 Vss 0.00410051f
c69 67 Vss 1.62518e-19
c70 62 Vss 7.10513e-22
c71 57 Vss 8.03422e-19
c72 52 Vss 9.77866e-19
c73 49 Vss 0.00537236f
c74 45 Vss 0.00387287f
c75 32 Vss 0.0350852f
c76 31 Vss 0.0994129f
c77 28 Vss 0.0350852f
c78 27 Vss 0.0994129f
c79 7 Vss 0.268864f
c80 3 Vss 0.268864f
r81 114 118 0.326018
r82 113 116 0.551426
r83 113 114 4.58464
r84 112 116 0.551426
r85 111 115 0.551426
r86 111 112 6.75193
r87 110 115 0.551426
r88 109 110 4.58464
r89 105 116 0.0828784
r90 101 115 0.0828784
r91 99 118 0.326018
r92 99 100 10.1279
r93 97 109 0.652036
r94 97 98 10.1279
r95 93 100 0.652036
r96 89 98 0.652036
r97 67 105 1.82344
r98 62 101 1.82344
r99 57 77 1.16709
r100 57 93 2.16729
r101 52 72 1.16709
r102 52 89 2.16729
r103 49 67 1.16709
r104 45 62 1.16709
r105 34 77 0.0476429
r106 32 34 1.45875
r107 31 38 0.652036
r108 31 34 1.45875
r109 30 72 0.0476429
r110 28 30 1.45875
r111 27 35 0.652036
r112 27 30 1.45875
r113 24 32 0.652036
r114 21 28 0.652036
r115 12 49 0.185659
r116 10 45 0.185659
r117 7 38 3.8511
r118 7 24 3.8511
r119 3 35 3.8511
r120 3 21 3.8511
.ends

.subckt PM_G2_BUF1_N2_A 2 4 12 22 28 Vss
c16 28 Vss 0.00294568f
c17 22 Vss 4.01518e-19
c18 12 Vss 0.200588f
c19 9 Vss 0.126125f
c20 7 Vss 0.0247918f
c21 4 Vss 0.139046f
r22 25 28 1.16709
r23 22 25 0.0416786
r24 15 28 0.0476429
r25 13 15 0.326018
r26 13 15 0.1167
r27 12 16 0.652036
r28 12 15 6.7686
r29 9 28 0.357321
r30 7 15 0.326018
r31 7 9 0.40845
r32 4 16 3.8511
r33 2 9 3.44265
.ends

.subckt PM_G2_BUF1_N2_Z 2 4 13 18 Vss
c14 18 Vss 4.84617e-19
c15 13 Vss 0.00522706f
c16 4 Vss 0.00176567f
r17 13 18 1.16709
r18 4 13 0.185659
r19 2 13 0.185659
.ends

.subckt PM_G2_BUF1_N2_NET17 2 4 6 8 18 33 36 41 50 58 Vss
c37 58 Vss 6.57973e-19
c38 50 Vss 0.00325633f
c39 41 Vss 0.00142824f
c40 36 Vss 0.00169654f
c41 33 Vss 0.00522706f
c42 22 Vss 0.0247918f
c43 19 Vss 0.0299669f
c44 18 Vss 0.169609f
c45 8 Vss 0.00176567f
c46 6 Vss 0.126125f
c47 2 Vss 0.138383f
r48 54 58 0.653045
r49 41 50 1.16709
r50 41 58 2.1395
r51 36 54 4.37625
r52 33 36 1.16709
r53 28 50 0.0476429
r54 26 50 0.357321
r55 22 28 0.326018
r56 22 26 0.40845
r57 19 28 6.7686
r58 18 28 0.326018
r59 18 28 0.1167
r60 15 19 0.652036
r61 8 33 0.185659
r62 6 26 3.44265
r63 4 33 0.185659
r64 2 15 3.8511
.ends

.subckt G2_BUF1_N2  VDD VSS A Z
*
* Z	Z
* A	A
* VSS	VSS
* VDD	VDD
XI10.X0 N_Z_XI10.X0_D N_VSS_XI10.X0_PGD N_NET17_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW8
XI7.X0 N_NET17_XI7.X0_D N_VSS_XI7.X0_PGD N_A_XI7.X0_CG N_VSS_XI7.X0_PGD
+ N_VDD_XI7.X0_S TIGFET_HPNW8
XI9.X0 N_Z_XI9.X0_D N_VDD_XI9.X0_PGD N_NET17_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW8
XI8.X0 N_NET17_XI8.X0_D N_VDD_XI8.X0_PGD N_A_XI8.X0_CG N_VDD_XI8.X0_PGD
+ N_VSS_XI8.X0_S TIGFET_HPNW8
*
x_PM_G2_BUF1_N2_VDD N_VDD_XI10.X0_S N_VDD_XI7.X0_S N_VDD_XI9.X0_PGD
+ N_VDD_XI8.X0_PGD N_VDD_c_4_p N_VDD_c_50_p N_VDD_c_8_p N_VDD_c_36_p
+ N_VDD_c_45_p N_VDD_c_6_p N_VDD_c_34_p N_VDD_c_3_p N_VDD_c_5_p N_VDD_c_38_p
+ N_VDD_c_46_p N_VDD_c_9_p N_VDD_c_13_p N_VDD_c_17_p VDD N_VDD_c_14_p
+ N_VDD_c_18_p Vss PM_G2_BUF1_N2_VDD
x_PM_G2_BUF1_N2_VSS N_VSS_XI10.X0_PGD N_VSS_XI7.X0_PGD N_VSS_XI9.X0_S
+ N_VSS_XI8.X0_S N_VSS_c_63_n N_VSS_c_65_n N_VSS_c_93_p N_VSS_c_67_n
+ N_VSS_c_69_n N_VSS_c_100_p N_VSS_c_106_p N_VSS_c_70_n N_VSS_c_74_n
+ N_VSS_c_101_p N_VSS_c_107_p N_VSS_c_78_n N_VSS_c_82_n N_VSS_c_85_n
+ N_VSS_c_86_n N_VSS_c_87_n N_VSS_c_88_n N_VSS_c_103_p N_VSS_c_110_p
+ N_VSS_c_89_n N_VSS_c_111_p N_VSS_c_90_n VSS Vss PM_G2_BUF1_N2_VSS
x_PM_G2_BUF1_N2_A N_A_XI7.X0_CG N_A_XI8.X0_CG N_A_c_116_n A N_A_c_119_n Vss
+ PM_G2_BUF1_N2_A
x_PM_G2_BUF1_N2_Z N_Z_XI10.X0_D N_Z_XI9.X0_D N_Z_c_132_n Z Vss PM_G2_BUF1_N2_Z
x_PM_G2_BUF1_N2_NET17 N_NET17_XI10.X0_CG N_NET17_XI7.X0_D N_NET17_XI9.X0_CG
+ N_NET17_XI8.X0_D N_NET17_c_147_n N_NET17_c_149_n N_NET17_c_151_n
+ N_NET17_c_154_n N_NET17_c_160_n N_NET17_c_163_n Vss PM_G2_BUF1_N2_NET17
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI10.X0_PGD 0.00201245f
cc_2 N_VDD_XI8.X0_PGD N_VSS_XI7.X0_PGD 0.00201245f
cc_3 N_VDD_c_3_p N_VSS_XI7.X0_PGD 3.05236e-19
cc_4 N_VDD_c_4_p N_VSS_c_63_n 0.00201245f
cc_5 N_VDD_c_5_p N_VSS_c_63_n 3.9313e-19
cc_6 N_VDD_c_6_p N_VSS_c_65_n 3.05236e-19
cc_7 N_VDD_c_5_p N_VSS_c_65_n 4.1253e-19
cc_8 N_VDD_c_8_p N_VSS_c_67_n 0.00201245f
cc_9 N_VDD_c_9_p N_VSS_c_67_n 3.9313e-19
cc_10 N_VDD_c_9_p N_VSS_c_69_n 4.1253e-19
cc_11 N_VDD_c_6_p N_VSS_c_70_n 8.67538e-19
cc_12 N_VDD_c_5_p N_VSS_c_70_n 0.00161703f
cc_13 N_VDD_c_13_p N_VSS_c_70_n 0.00106273f
cc_14 N_VDD_c_14_p N_VSS_c_70_n 3.48267e-19
cc_15 N_VDD_c_3_p N_VSS_c_74_n 8.67538e-19
cc_16 N_VDD_c_9_p N_VSS_c_74_n 0.00161703f
cc_17 N_VDD_c_17_p N_VSS_c_74_n 0.00110056f
cc_18 N_VDD_c_18_p N_VSS_c_74_n 3.48267e-19
cc_19 N_VDD_c_6_p N_VSS_c_78_n 3.66936e-19
cc_20 N_VDD_c_5_p N_VSS_c_78_n 2.26455e-19
cc_21 N_VDD_c_13_p N_VSS_c_78_n 3.99794e-19
cc_22 N_VDD_c_14_p N_VSS_c_78_n 6.489e-19
cc_23 N_VDD_c_3_p N_VSS_c_82_n 3.66936e-19
cc_24 N_VDD_c_9_p N_VSS_c_82_n 2.26455e-19
cc_25 N_VDD_c_18_p N_VSS_c_82_n 6.489e-19
cc_26 N_VDD_c_5_p N_VSS_c_85_n 0.00567457f
cc_27 N_VDD_c_5_p N_VSS_c_86_n 0.0017359f
cc_28 N_VDD_c_9_p N_VSS_c_87_n 0.00573644f
cc_29 N_VDD_c_9_p N_VSS_c_88_n 0.0017359f
cc_30 N_VDD_c_13_p N_VSS_c_89_n 3.85245e-19
cc_31 N_VDD_c_17_p N_VSS_c_90_n 3.85245e-19
cc_32 N_VDD_XI9.X0_PGD N_A_c_116_n 4.12647e-19
cc_33 N_VDD_XI8.X0_PGD N_A_c_116_n 4.07423e-19
cc_34 N_VDD_c_34_p A 9.3432e-19
cc_35 N_VDD_c_34_p N_A_c_119_n 5.18354e-19
cc_36 N_VDD_c_36_p N_Z_c_132_n 3.43419e-19
cc_37 N_VDD_c_5_p N_Z_c_132_n 3.4118e-19
cc_38 N_VDD_c_38_p N_Z_c_132_n 3.72199e-19
cc_39 N_VDD_c_36_p Z 3.48267e-19
cc_40 N_VDD_c_5_p Z 4.58391e-19
cc_41 N_VDD_c_38_p Z 7.4527e-19
cc_42 N_VDD_c_34_p N_NET17_XI10.X0_CG 2.86271e-19
cc_43 N_VDD_XI9.X0_PGD N_NET17_c_147_n 4.07423e-19
cc_44 N_VDD_XI8.X0_PGD N_NET17_c_147_n 4.12647e-19
cc_45 N_VDD_c_45_p N_NET17_c_149_n 3.43419e-19
cc_46 N_VDD_c_46_p N_NET17_c_149_n 3.72199e-19
cc_47 N_VDD_c_45_p N_NET17_c_151_n 3.48267e-19
cc_48 N_VDD_c_46_p N_NET17_c_151_n 8.0086e-19
cc_49 N_VDD_c_9_p N_NET17_c_151_n 4.34701e-19
cc_50 N_VDD_c_50_p N_NET17_c_154_n 3.02565e-19
cc_51 N_VDD_c_34_p N_NET17_c_154_n 2.74452e-19
cc_52 N_VDD_c_13_p N_NET17_c_154_n 4.44912e-19
cc_53 N_VDD_c_17_p N_NET17_c_154_n 2.83214e-19
cc_54 N_VDD_c_14_p N_NET17_c_154_n 3.49905e-19
cc_55 N_VDD_c_18_p N_NET17_c_154_n 4.45791e-19
cc_56 N_VDD_c_13_p N_NET17_c_160_n 3.43988e-19
cc_57 N_VDD_c_17_p N_NET17_c_160_n 2.24759e-19
cc_58 N_VDD_c_14_p N_NET17_c_160_n 2.68747e-19
cc_59 N_VDD_c_34_p N_NET17_c_163_n 4.34465e-19
cc_60 N_VSS_XI10.X0_PGD N_A_c_116_n 4.12647e-19
cc_61 N_VSS_XI7.X0_PGD N_A_c_116_n 4.04227e-19
cc_62 N_VSS_c_93_p A 2.23478e-19
cc_63 N_VSS_c_74_n A 3.28992e-19
cc_64 N_VSS_c_78_n A 2.26741e-19
cc_65 N_VSS_c_82_n A 6.58807e-19
cc_66 N_VSS_c_70_n N_A_c_119_n 2.11378e-19
cc_67 N_VSS_c_74_n N_A_c_119_n 3.2351e-19
cc_68 N_VSS_c_82_n N_A_c_119_n 2.68747e-19
cc_69 N_VSS_c_100_p N_Z_c_132_n 3.43419e-19
cc_70 N_VSS_c_101_p N_Z_c_132_n 3.48267e-19
cc_71 N_VSS_c_101_p Z 5.37696e-19
cc_72 N_VSS_c_103_p Z 2.7826e-19
cc_73 N_VSS_XI10.X0_PGD N_NET17_c_147_n 4.04227e-19
cc_74 N_VSS_XI7.X0_PGD N_NET17_c_147_n 4.12647e-19
cc_75 N_VSS_c_106_p N_NET17_c_149_n 3.43419e-19
cc_76 N_VSS_c_107_p N_NET17_c_149_n 3.48267e-19
cc_77 N_VSS_c_107_p N_NET17_c_151_n 4.8288e-19
cc_78 N_VSS_c_87_n N_NET17_c_151_n 4.84973e-19
cc_79 N_VSS_c_110_p N_NET17_c_151_n 5.49885e-19
cc_80 N_VSS_c_111_p N_NET17_c_151_n 0.00103514f
cc_81 N_VSS_c_85_n N_NET17_c_154_n 2.50699e-19
cc_82 N_VSS_c_111_p N_NET17_c_154_n 0.00119345f
cc_83 N_VSS_c_85_n N_NET17_c_163_n 8.43205e-19
cc_84 N_VSS_c_87_n N_NET17_c_163_n 4.88529e-19
cc_85 N_A_c_116_n N_NET17_c_147_n 0.0093393f
cc_86 N_A_c_116_n N_NET17_c_149_n 4.95639e-19
cc_87 A N_NET17_c_151_n 8.54729e-19
cc_88 N_Z_c_132_n N_NET17_c_147_n 4.95639e-19
cc_89 N_Z_c_132_n N_NET17_c_149_n 4.64289e-19
cc_90 Z N_NET17_c_149_n 2.11378e-19
cc_91 N_Z_c_132_n N_NET17_c_151_n 2.11378e-19
*
.ends
*
*
.subckt BUF1_HPNW8 A Y VDD VSS
xgate (VDD VSS A Y) G2_BUF1_N2
.ends
*
* File: G3_DFFQ1_N2.pex.netlist
* Created: Wed Apr  6 11:10:43 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_DFFQ1_N2_VSS 2 4 6 8 10 12 14 29 42 44 49 55 59 64 67 72 78 83 88
+ 93 102 111 116 125 126 127 128 132 137 142 148 154 156 161 163 165 166 167 Vss
c103 167 Vss 4.28045e-19
c104 166 Vss 3.75522e-19
c105 165 Vss 3.75522e-19
c106 164 Vss 6.15603e-19
c107 163 Vss 0.00495722f
c108 161 Vss 0.0016477f
c109 156 Vss 0.00136752f
c110 154 Vss 0.00253212f
c111 148 Vss 0.004602f
c112 142 Vss 0.00300844f
c113 132 Vss 0.0019674f
c114 128 Vss 6.73974e-19
c115 127 Vss 8.13835e-19
c116 126 Vss 0.00570183f
c117 125 Vss 0.00160501f
c118 116 Vss 0.00497548f
c119 111 Vss 0.00376876f
c120 102 Vss 0.00442938f
c121 93 Vss 2.73987e-19
c122 88 Vss 8.09754e-19
c123 83 Vss 7.28045e-19
c124 78 Vss 0.00155391f
c125 72 Vss 0.0108629f
c126 67 Vss 0.00135556f
c127 64 Vss 0.00650697f
c128 59 Vss 0.00498022f
c129 55 Vss 0.00373197f
c130 49 Vss 0.0568987f
c131 44 Vss 0.0568992f
c132 42 Vss 1.04992e-19
c133 29 Vss 0.035607f
c134 28 Vss 0.101294f
c135 14 Vss 0.134651f
c136 8 Vss 0.136772f
c137 6 Vss 0.133795f
c138 4 Vss 0.133902f
r139 162 167 0.551426
r140 162 163 15.5878
r141 161 167 0.551426
r142 160 161 4.62632
r143 156 167 0.0828784
r144 155 166 0.494161
r145 154 163 0.652036
r146 154 155 4.37625
r147 150 166 0.128424
r148 149 165 0.494161
r149 148 160 0.652036
r150 148 149 10.1279
r151 144 165 0.128424
r152 143 164 0.494161
r153 142 166 0.494161
r154 142 143 7.46046
r155 138 164 0.128424
r156 132 164 0.494161
r157 132 137 1.00029
r158 126 165 0.494161
r159 126 127 15.8795
r160 125 128 0.655813
r161 124 127 0.652036
r162 124 125 4.62632
r163 93 156 1.82344
r164 88 116 1.16709
r165 88 150 2.16729
r166 83 111 1.16709
r167 83 144 2.16729
r168 78 138 5.2515
r169 75 137 1.29204
r170 72 102 1.16709
r171 72 75 13.7539
r172 67 128 1.82344
r173 64 93 1.16709
r174 59 78 1.16709
r175 55 67 1.16709
r176 49 116 0.197068
r177 46 49 1.2837
r178 42 111 0.197068
r179 42 44 1.2837
r180 38 46 0.0685365
r181 35 44 0.0685365
r182 31 102 0.0476429
r183 29 31 1.45875
r184 28 32 0.652036
r185 28 31 1.45875
r186 25 29 0.652036
r187 14 38 3.8511
r188 12 64 0.185659
r189 10 59 0.185659
r190 8 35 3.8511
r191 6 32 3.8511
r192 4 25 3.8511
r193 2 55 0.185659
.ends

.subckt PM_G3_DFFQ1_N2_CK 2 4 6 8 18 21 25 37 40 Vss
c33 40 Vss 0.00476958f
c34 37 Vss 3.41336e-19
c35 33 Vss 0.0299314f
c36 25 Vss 0.166342f
c37 21 Vss 1.04992e-19
c38 18 Vss 0.18663f
c39 15 Vss 0.12596f
c40 13 Vss 0.0247918f
c41 6 Vss 0.550304f
c42 4 Vss 0.136627f
r43 37 40 1.16709
r44 26 33 0.494161
r45 25 27 0.652036
r46 25 26 4.84305
r47 22 33 0.128424
r48 21 40 0.0238214
r49 19 21 0.326018
r50 19 21 0.1167
r51 18 33 0.494161
r52 18 21 6.7686
r53 15 40 0.357321
r54 13 21 0.326018
r55 13 15 0.3501
r56 6 8 15.4044
r57 6 27 3.8511
r58 4 22 3.8511
r59 2 15 3.501
.ends

.subckt PM_G3_DFFQ1_N2_VDD 2 4 6 8 10 12 14 28 42 44 49 56 60 63 64 65 70 72 76
+ 78 79 82 84 86 91 93 95 96 98 99 100 102 104 113 118 Vss
c109 118 Vss 0.00535583f
c110 113 Vss 0.00546246f
c111 104 Vss 0.00475709f
c112 100 Vss 4.52364e-19
c113 99 Vss 2.39889e-19
c114 98 Vss 4.42806e-19
c115 96 Vss 0.00368915f
c116 95 Vss 5.05789e-19
c117 93 Vss 0.00304576f
c118 91 Vss 0.00856613f
c119 86 Vss 0.00179444f
c120 84 Vss 0.00304688f
c121 82 Vss 0.00102756f
c122 79 Vss 4.90412e-19
c123 78 Vss 0.00536329f
c124 76 Vss 6.6871e-19
c125 72 Vss 0.00341969f
c126 70 Vss 0.00232792f
c127 67 Vss 0.00182492f
c128 65 Vss 8.64465e-19
c129 64 Vss 0.00774944f
c130 63 Vss 0.00502551f
c131 60 Vss 0.00655192f
c132 56 Vss 0.00779243f
c133 49 Vss 0.0588939f
c134 44 Vss 0.0581359f
c135 42 Vss 1.01357e-19
c136 29 Vss 0.0372896f
c137 28 Vss 0.10099f
c138 12 Vss 0.13719f
c139 10 Vss 0.13484f
c140 8 Vss 0.00143442f
c141 4 Vss 0.136142f
c142 2 Vss 0.134971f
r143 95 104 1.16709
r144 95 96 0.470345
r145 93 102 0.326018
r146 92 100 0.551426
r147 92 93 4.58464
r148 91 100 0.551426
r149 90 91 15.6295
r150 86 100 0.0828784
r151 86 88 1.82344
r152 85 99 0.494161
r153 84 90 0.652036
r154 84 85 4.37625
r155 82 118 1.16709
r156 80 99 0.128424
r157 80 82 2.16729
r158 78 102 0.326018
r159 78 79 10.1279
r160 76 113 1.16709
r161 74 79 0.652036
r162 74 76 2.16729
r163 73 98 0.494161
r164 72 99 0.494161
r165 72 73 7.46046
r166 68 98 0.128424
r167 68 70 5.29318
r168 67 96 3.82922
r169 64 98 0.494161
r170 64 65 13.0037
r171 63 67 0.655813
r172 62 65 0.652036
r173 62 63 8.37739
r174 60 88 1.16709
r175 56 70 1.16709
r176 49 118 0.197068
r177 46 49 1.2837
r178 42 113 0.197068
r179 42 44 1.2837
r180 38 46 0.0685365
r181 35 44 0.0685365
r182 31 104 0.0476429
r183 29 31 1.45875
r184 28 32 0.652036
r185 28 31 1.45875
r186 25 29 0.652036
r187 14 60 0.185659
r188 12 38 3.8511
r189 10 35 3.8511
r190 8 56 0.185659
r191 6 56 0.185659
r192 4 25 3.8511
r193 2 32 3.8511
.ends

.subckt PM_G3_DFFQ1_N2_CKN 2 4 6 8 18 25 28 33 50 Vss
c38 51 Vss 0.00128326f
c39 50 Vss 0.00576518f
c40 33 Vss 7.37543e-19
c41 28 Vss 0.00177951f
c42 25 Vss 0.00542517f
c43 18 Vss 7.82969e-19
c44 6 Vss 0.475302f
c45 4 Vss 0.00143442f
r46 50 51 14.6709
r47 46 51 0.652036
r48 33 50 0.531835
r49 28 46 4.91807
r50 25 28 1.16709
r51 18 33 1.16709
r52 8 18 7.7022
r53 6 18 7.7022
r54 4 25 0.185659
r55 2 25 0.185659
.ends

.subckt PM_G3_DFFQ1_N2_D 2 4 11 12 22 25 28 Vss
c24 28 Vss 0.00170116f
c25 25 Vss 4.81931e-19
c26 12 Vss 0.21156f
c27 11 Vss 9.81474e-20
c28 7 Vss 0.0247918f
c29 4 Vss 0.137342f
c30 2 Vss 0.125849f
r31 25 28 1.16709
r32 22 25 0.0364688
r33 15 28 0.0476429
r34 13 15 0.326018
r35 13 15 0.1167
r36 12 16 0.652036
r37 12 15 6.7686
r38 11 28 0.357321
r39 7 15 0.326018
r40 7 11 0.40845
r41 4 16 3.8511
r42 2 11 3.44265
.ends

.subckt PM_G3_DFFQ1_N2_X 2 4 6 8 17 20 23 33 35 39 41 47 Vss
c47 47 Vss 0.00138877f
c48 41 Vss 5.3862e-19
c49 39 Vss 0.00123905f
c50 35 Vss 0.00217266f
c51 33 Vss 0.00551754f
c52 23 Vss 1.01432e-19
c53 20 Vss 0.21178f
c54 17 Vss 0.125802f
c55 15 Vss 0.0247918f
c56 8 Vss 0.137267f
c57 6 Vss 0.00143442f
r58 44 47 1.16709
r59 41 44 2.08393
r60 37 39 5.2515
r61 36 41 0.0685365
r62 35 37 0.652036
r63 35 36 1.70882
r64 33 39 1.16709
r65 23 47 0.0476429
r66 21 23 0.326018
r67 21 23 0.1167
r68 20 24 0.652036
r69 20 23 6.7686
r70 17 47 0.357321
r71 15 23 0.326018
r72 15 17 0.40845
r73 8 24 3.8511
r74 6 33 0.185659
r75 4 17 3.44265
r76 2 33 0.185659
.ends

.subckt PM_G3_DFFQ1_N2_Q 2 4 13 16 Vss
c12 16 Vss 3.81501e-19
c13 13 Vss 0.00450389f
c14 4 Vss 0.00143442f
r15 16 19 0.0416786
r16 13 19 1.16709
r17 4 13 0.185659
r18 2 13 0.185659
.ends

.subckt G3_DFFQ1_N2  VSS CK VDD D Q
*
* Q	Q
* D	D
* VDD	VDD
* CK	CK
* VSS	VSS
XI6.X0 N_CKN_XI6.X0_D N_VDD_XI6.X0_PGD N_CK_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW8
XI7.X0 N_CKN_XI7.X0_D N_VSS_XI7.X0_PGD N_CK_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW8
XI11.X0 N_X_XI11.X0_D N_VSS_XI11.X0_PGD N_D_XI11.X0_CG N_CK_XI11.X0_PGS
+ N_VDD_XI11.X0_S TIGFET_HPNW8
XI8.X0 N_Q_XI8.X0_D N_VDD_XI8.X0_PGD N_X_XI8.X0_CG N_CK_XI8.X0_PGS
+ N_VSS_XI8.X0_S TIGFET_HPNW8
XI10.X0 N_X_XI10.X0_D N_VDD_XI10.X0_PGD N_D_XI10.X0_CG N_CKN_XI10.X0_PGS
+ N_VSS_XI10.X0_S TIGFET_HPNW8
XI9.X0 N_Q_XI9.X0_D N_VSS_XI9.X0_PGD N_X_XI9.X0_CG N_CKN_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW8
*
x_PM_G3_DFFQ1_N2_VSS N_VSS_XI6.X0_S N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS
+ N_VSS_XI11.X0_PGD N_VSS_XI8.X0_S N_VSS_XI10.X0_S N_VSS_XI9.X0_PGD N_VSS_c_11_p
+ N_VSS_c_80_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_14_p N_VSS_c_101_p N_VSS_c_91_p
+ N_VSS_c_15_p N_VSS_c_3_p N_VSS_c_30_p N_VSS_c_21_p N_VSS_c_31_p N_VSS_c_41_p
+ N_VSS_c_53_p N_VSS_c_4_p N_VSS_c_34_p N_VSS_c_16_p N_VSS_c_7_p N_VSS_c_20_p
+ N_VSS_c_17_p N_VSS_c_77_p VSS N_VSS_c_35_p N_VSS_c_27_p N_VSS_c_36_p
+ N_VSS_c_43_p N_VSS_c_45_p N_VSS_c_46_p N_VSS_c_28_p N_VSS_c_37_p N_VSS_c_47_p
+ Vss PM_G3_DFFQ1_N2_VSS
x_PM_G3_DFFQ1_N2_CK N_CK_XI6.X0_CG N_CK_XI7.X0_CG N_CK_XI11.X0_PGS
+ N_CK_XI8.X0_PGS N_CK_c_108_n N_CK_c_125_p N_CK_c_109_n CK N_CK_c_115_p Vss
+ PM_G3_DFFQ1_N2_CK
x_PM_G3_DFFQ1_N2_VDD N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI7.X0_S
+ N_VDD_XI11.X0_S N_VDD_XI8.X0_PGD N_VDD_XI10.X0_PGD N_VDD_XI9.X0_S
+ N_VDD_c_140_n N_VDD_c_227_p N_VDD_c_141_n N_VDD_c_142_n N_VDD_c_214_p
+ N_VDD_c_240_p N_VDD_c_143_n N_VDD_c_147_n N_VDD_c_149_n N_VDD_c_150_n
+ N_VDD_c_152_n N_VDD_c_158_n N_VDD_c_161_n N_VDD_c_167_n N_VDD_c_168_n
+ N_VDD_c_170_n N_VDD_c_172_n N_VDD_c_173_n N_VDD_c_177_n N_VDD_c_181_n
+ N_VDD_c_183_n N_VDD_c_185_n N_VDD_c_186_n N_VDD_c_187_n VDD N_VDD_c_188_n
+ N_VDD_c_190_n N_VDD_c_193_n Vss PM_G3_DFFQ1_N2_VDD
x_PM_G3_DFFQ1_N2_CKN N_CKN_XI6.X0_D N_CKN_XI7.X0_D N_CKN_XI10.X0_PGS
+ N_CKN_XI9.X0_PGS N_CKN_c_261_n N_CKN_c_246_n N_CKN_c_248_n N_CKN_c_252_n
+ N_CKN_c_253_n Vss PM_G3_DFFQ1_N2_CKN
x_PM_G3_DFFQ1_N2_D N_D_XI11.X0_CG N_D_XI10.X0_CG N_D_c_284_n N_D_c_285_n D
+ N_D_c_286_n N_D_c_290_n Vss PM_G3_DFFQ1_N2_D
x_PM_G3_DFFQ1_N2_X N_X_XI11.X0_D N_X_XI8.X0_CG N_X_XI10.X0_D N_X_XI9.X0_CG
+ N_X_c_320_n N_X_c_308_n N_X_c_323_n N_X_c_309_n N_X_c_311_n N_X_c_312_n
+ N_X_c_316_n N_X_c_318_n Vss PM_G3_DFFQ1_N2_X
x_PM_G3_DFFQ1_N2_Q N_Q_XI8.X0_D N_Q_XI9.X0_D N_Q_c_355_n Q Vss PM_G3_DFFQ1_N2_Q
cc_1 N_VSS_XI7.X0_PGS N_CK_XI11.X0_PGS 0.00316278f
cc_2 N_VSS_XI11.X0_PGD N_CK_XI11.X0_PGS 0.00164185f
cc_3 N_VSS_c_3_p N_CK_XI11.X0_PGS 8.34822e-19
cc_4 N_VSS_c_4_p N_CK_XI11.X0_PGS 4.02129e-19
cc_5 N_VSS_XI7.X0_PGD N_CK_c_108_n 4.18808e-19
cc_6 N_VSS_XI7.X0_PGS N_CK_c_109_n 4.29708e-19
cc_7 N_VSS_c_7_p CK 5.33707e-19
cc_8 N_VSS_XI7.X0_PGD N_VDD_XI6.X0_PGD 0.00196344f
cc_9 N_VSS_XI9.X0_PGD N_VDD_XI8.X0_PGD 0.00221773f
cc_10 N_VSS_XI11.X0_PGD N_VDD_XI10.X0_PGD 0.00211593f
cc_11 N_VSS_c_11_p N_VDD_c_140_n 0.00196344f
cc_12 N_VSS_c_12_p N_VDD_c_141_n 0.00221773f
cc_13 N_VSS_c_13_p N_VDD_c_142_n 0.00211593f
cc_14 N_VSS_c_14_p N_VDD_c_143_n 9.5668e-19
cc_15 N_VSS_c_15_p N_VDD_c_143_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_143_n 0.00352032f
cc_17 N_VSS_c_17_p N_VDD_c_143_n 0.00185572f
cc_18 N_VSS_c_15_p N_VDD_c_147_n 4.50735e-19
cc_19 N_VSS_c_7_p N_VDD_c_147_n 0.00936712f
cc_20 N_VSS_c_20_p N_VDD_c_149_n 0.00105561f
cc_21 N_VSS_c_21_p N_VDD_c_150_n 0.00233232f
cc_22 N_VSS_c_4_p N_VDD_c_150_n 9.47758e-19
cc_23 N_VSS_c_13_p N_VDD_c_152_n 2.74851e-19
cc_24 N_VSS_c_21_p N_VDD_c_152_n 0.00161703f
cc_25 N_VSS_c_4_p N_VDD_c_152_n 2.24973e-19
cc_26 N_VSS_c_7_p N_VDD_c_152_n 0.00133545f
cc_27 N_VSS_c_27_p N_VDD_c_152_n 0.00408783f
cc_28 N_VSS_c_28_p N_VDD_c_152_n 7.74609e-19
cc_29 N_VSS_c_3_p N_VDD_c_158_n 0.00179097f
cc_30 N_VSS_c_30_p N_VDD_c_158_n 3.92901e-19
cc_31 N_VSS_c_31_p N_VDD_c_158_n 8.83788e-19
cc_32 N_VSS_c_12_p N_VDD_c_161_n 3.66315e-19
cc_33 N_VSS_c_31_p N_VDD_c_161_n 0.00141228f
cc_34 N_VSS_c_34_p N_VDD_c_161_n 0.00114511f
cc_35 N_VSS_c_35_p N_VDD_c_161_n 0.00409335f
cc_36 N_VSS_c_36_p N_VDD_c_161_n 0.00330569f
cc_37 N_VSS_c_37_p N_VDD_c_161_n 7.74609e-19
cc_38 N_VSS_c_35_p N_VDD_c_167_n 0.00144699f
cc_39 N_VSS_c_21_p N_VDD_c_168_n 9.29349e-19
cc_40 N_VSS_c_4_p N_VDD_c_168_n 3.79458e-19
cc_41 N_VSS_c_41_p N_VDD_c_170_n 4.50735e-19
cc_42 N_VSS_c_27_p N_VDD_c_170_n 0.00438429f
cc_43 N_VSS_c_43_p N_VDD_c_172_n 4.68065e-19
cc_44 N_VSS_c_41_p N_VDD_c_173_n 0.00187494f
cc_45 N_VSS_c_45_p N_VDD_c_173_n 0.00345634f
cc_46 N_VSS_c_46_p N_VDD_c_173_n 0.00778647f
cc_47 N_VSS_c_47_p N_VDD_c_173_n 9.16632e-19
cc_48 N_VSS_c_31_p N_VDD_c_177_n 4.35319e-19
cc_49 N_VSS_c_34_p N_VDD_c_177_n 3.66936e-19
cc_50 N_VSS_c_36_p N_VDD_c_177_n 0.00106857f
cc_51 N_VSS_c_46_p N_VDD_c_177_n 0.00335989f
cc_52 N_VSS_c_3_p N_VDD_c_181_n 6.19689e-19
cc_53 N_VSS_c_53_p N_VDD_c_181_n 3.8721e-19
cc_54 N_VSS_c_15_p N_VDD_c_183_n 0.00222015f
cc_55 N_VSS_c_7_p N_VDD_c_183_n 2.66524e-19
cc_56 N_VSS_c_7_p N_VDD_c_185_n 0.00118128f
cc_57 N_VSS_c_27_p N_VDD_c_186_n 0.0010448f
cc_58 N_VSS_c_46_p N_VDD_c_187_n 0.00116512f
cc_59 N_VSS_c_3_p N_VDD_c_188_n 3.86162e-19
cc_60 N_VSS_c_53_p N_VDD_c_188_n 6.0892e-19
cc_61 N_VSS_c_3_p N_VDD_c_190_n 5.2607e-19
cc_62 N_VSS_c_31_p N_VDD_c_190_n 3.48267e-19
cc_63 N_VSS_c_34_p N_VDD_c_190_n 6.489e-19
cc_64 N_VSS_c_21_p N_VDD_c_193_n 3.48267e-19
cc_65 N_VSS_c_4_p N_VDD_c_193_n 6.20986e-19
cc_66 N_VSS_c_14_p N_CKN_c_246_n 3.43419e-19
cc_67 N_VSS_c_15_p N_CKN_c_246_n 3.48267e-19
cc_68 N_VSS_c_15_p N_CKN_c_248_n 0.00109746f
cc_69 N_VSS_c_3_p N_CKN_c_248_n 6.97825e-19
cc_70 N_VSS_c_7_p N_CKN_c_248_n 4.81255e-19
cc_71 N_VSS_c_46_p N_CKN_c_248_n 2.6973e-19
cc_72 N_VSS_c_46_p N_CKN_c_252_n 0.00111539f
cc_73 N_VSS_c_3_p N_CKN_c_253_n 0.00225294f
cc_74 N_VSS_c_30_p N_CKN_c_253_n 7.04847e-19
cc_75 N_VSS_c_31_p N_CKN_c_253_n 6.45464e-19
cc_76 N_VSS_c_7_p N_CKN_c_253_n 0.00132819f
cc_77 N_VSS_c_77_p N_CKN_c_253_n 7.24142e-19
cc_78 N_VSS_c_35_p N_CKN_c_253_n 7.58219e-19
cc_79 N_VSS_c_27_p N_CKN_c_253_n 9.23091e-19
cc_80 N_VSS_c_80_p N_D_c_284_n 9.24646e-19
cc_81 N_VSS_XI11.X0_PGD N_D_c_285_n 3.94389e-19
cc_82 N_VSS_c_3_p N_D_c_286_n 6.13924e-19
cc_83 N_VSS_c_21_p N_D_c_286_n 2.96367e-19
cc_84 N_VSS_c_53_p N_D_c_286_n 3.48267e-19
cc_85 N_VSS_c_4_p N_D_c_286_n 3.20302e-19
cc_86 N_VSS_c_3_p N_D_c_290_n 3.48267e-19
cc_87 N_VSS_c_21_p N_D_c_290_n 3.20302e-19
cc_88 N_VSS_c_53_p N_D_c_290_n 6.88619e-19
cc_89 N_VSS_c_4_p N_D_c_290_n 2.62417e-19
cc_90 N_VSS_XI9.X0_PGD N_X_c_308_n 4.04227e-19
cc_91 N_VSS_c_91_p N_X_c_309_n 3.43419e-19
cc_92 N_VSS_c_41_p N_X_c_309_n 3.48267e-19
cc_93 N_VSS_c_35_p N_X_c_311_n 2.44303e-19
cc_94 N_VSS_c_91_p N_X_c_312_n 3.48267e-19
cc_95 N_VSS_c_3_p N_X_c_312_n 4.71026e-19
cc_96 N_VSS_c_41_p N_X_c_312_n 5.71987e-19
cc_97 N_VSS_c_46_p N_X_c_312_n 2.97611e-19
cc_98 N_VSS_c_3_p N_X_c_316_n 0.00157847f
cc_99 N_VSS_c_46_p N_X_c_316_n 2.88807e-19
cc_100 N_VSS_c_3_p N_X_c_318_n 3.48267e-19
cc_101 N_VSS_c_101_p N_Q_c_355_n 3.43419e-19
cc_102 N_VSS_c_30_p N_Q_c_355_n 3.48267e-19
cc_103 N_VSS_c_30_p Q 5.37696e-19
cc_104 N_CK_c_108_n N_VDD_XI6.X0_PGD 4.18808e-19
cc_105 N_CK_XI11.X0_PGS N_VDD_XI10.X0_PGD 2.44781e-19
cc_106 N_CK_c_109_n N_VDD_c_142_n 2.44781e-19
cc_107 CK N_VDD_c_143_n 5.04211e-19
cc_108 N_CK_c_115_p N_VDD_c_143_n 5.30123e-19
cc_109 N_CK_c_108_n N_VDD_c_147_n 0.0015171f
cc_110 CK N_VDD_c_147_n 0.00141439f
cc_111 N_CK_c_115_p N_VDD_c_147_n 0.00120239f
cc_112 N_CK_XI11.X0_PGS N_VDD_c_150_n 2.48209e-19
cc_113 N_CK_c_109_n N_VDD_c_150_n 5.56076e-19
cc_114 CK N_VDD_c_150_n 3.85155e-19
cc_115 N_CK_c_115_p N_VDD_c_150_n 2.72301e-19
cc_116 CK N_VDD_c_181_n 4.2144e-19
cc_117 N_CK_c_115_p N_VDD_c_181_n 3.27641e-19
cc_118 N_CK_c_125_p N_VDD_c_188_n 9.40274e-19
cc_119 CK N_VDD_c_188_n 3.20302e-19
cc_120 N_CK_c_115_p N_VDD_c_188_n 2.62417e-19
cc_121 N_CK_XI11.X0_PGS N_CKN_XI10.X0_PGS 4.11563e-19
cc_122 N_CK_XI11.X0_PGS N_CKN_c_261_n 2.73384e-19
cc_123 N_CK_c_108_n N_CKN_c_246_n 6.55689e-19
cc_124 N_CK_XI11.X0_PGS N_D_XI11.X0_CG 4.28946e-19
cc_125 N_CK_XI11.X0_PGS N_D_XI10.X0_CG 2.59344e-19
cc_126 N_CK_XI11.X0_PGS N_D_c_290_n 0.00300565f
cc_127 N_CK_XI11.X0_PGS N_X_XI9.X0_CG 2.61247e-19
cc_128 N_CK_XI11.X0_PGS N_X_c_320_n 4.55333e-19
cc_129 N_CK_XI11.X0_PGS N_X_c_318_n 0.00630896f
cc_130 N_VDD_c_173_n N_CKN_XI10.X0_PGS 7.25969e-19
cc_131 N_VDD_c_173_n N_CKN_c_261_n 8.21431e-19
cc_132 N_VDD_c_214_p N_CKN_c_246_n 3.43419e-19
cc_133 N_VDD_c_214_p N_CKN_c_248_n 3.48267e-19
cc_134 N_VDD_c_143_n N_CKN_c_248_n 3.84058e-19
cc_135 N_VDD_c_147_n N_CKN_c_248_n 4.28606e-19
cc_136 N_VDD_c_150_n N_CKN_c_248_n 5.37696e-19
cc_137 N_VDD_c_181_n N_CKN_c_248_n 6.42405e-19
cc_138 N_VDD_c_173_n N_CKN_c_252_n 7.71262e-19
cc_139 N_VDD_c_147_n N_CKN_c_253_n 3.98085e-19
cc_140 N_VDD_c_152_n N_CKN_c_253_n 2.80228e-19
cc_141 N_VDD_c_161_n N_CKN_c_253_n 4.0976e-19
cc_142 N_VDD_c_168_n N_CKN_c_253_n 2.45963e-19
cc_143 N_VDD_XI10.X0_PGD N_D_c_285_n 4.07433e-19
cc_144 N_VDD_XI8.X0_PGD N_X_c_308_n 3.96342e-19
cc_145 N_VDD_c_227_p N_X_c_323_n 8.75838e-19
cc_146 N_VDD_c_214_p N_X_c_309_n 3.43419e-19
cc_147 N_VDD_c_150_n N_X_c_309_n 3.48267e-19
cc_148 N_VDD_c_152_n N_X_c_309_n 3.37713e-19
cc_149 N_VDD_c_214_p N_X_c_312_n 3.48267e-19
cc_150 N_VDD_c_150_n N_X_c_312_n 6.94315e-19
cc_151 N_VDD_c_152_n N_X_c_312_n 4.72817e-19
cc_152 N_VDD_c_173_n N_X_c_312_n 0.00111552f
cc_153 N_VDD_c_158_n N_X_c_316_n 4.35824e-19
cc_154 N_VDD_c_173_n N_X_c_316_n 2.02855e-19
cc_155 N_VDD_c_190_n N_X_c_316_n 3.40502e-19
cc_156 N_VDD_c_158_n N_X_c_318_n 3.43988e-19
cc_157 N_VDD_c_190_n N_X_c_318_n 2.68747e-19
cc_158 N_VDD_c_240_p N_Q_c_355_n 3.43419e-19
cc_159 N_VDD_c_161_n N_Q_c_355_n 3.4118e-19
cc_160 N_VDD_c_172_n N_Q_c_355_n 3.72199e-19
cc_161 N_VDD_c_240_p Q 3.48267e-19
cc_162 N_VDD_c_161_n Q 4.58391e-19
cc_163 N_VDD_c_172_n Q 7.06537e-19
cc_164 N_CKN_XI10.X0_PGS N_D_XI10.X0_CG 0.00419505f
cc_165 N_CKN_XI10.X0_PGS N_X_c_308_n 0.00425073f
cc_166 N_CKN_c_261_n N_X_c_311_n 5.71169e-19
cc_167 N_CKN_c_253_n N_X_c_311_n 0.00127072f
cc_168 N_CKN_c_248_n N_X_c_312_n 4.96487e-19
cc_169 N_CKN_c_252_n N_X_c_312_n 8.08281e-19
cc_170 N_CKN_c_253_n N_X_c_312_n 6.84099e-19
cc_171 N_CKN_c_253_n N_X_c_316_n 8.25313e-19
cc_172 N_D_c_285_n N_X_c_308_n 0.00474388f
cc_173 N_D_c_285_n N_X_c_309_n 6.8653e-19
cc_174 N_D_c_285_n N_X_c_312_n 3.40033e-19
cc_175 N_D_c_286_n N_X_c_312_n 0.00151909f
cc_176 N_D_c_290_n N_X_c_312_n 0.00104518f
cc_177 N_D_c_286_n N_X_c_316_n 0.00146206f
cc_178 N_D_c_290_n N_X_c_316_n 0.00103457f
cc_179 N_D_c_286_n N_X_c_318_n 4.56568e-19
cc_180 N_D_c_290_n N_X_c_318_n 0.00373359f
cc_181 N_X_c_308_n N_Q_c_355_n 6.8653e-19
cc_182 N_X_c_311_n N_Q_c_355_n 4.47287e-19
cc_183 N_X_c_311_n Q 6.7453e-19
*
.ends
*
*
.subckt DFFQ1_HPNW8 CK D Q VDD VSS
xgate (VSS CK VDD D Q) G3_DFFQ1_N2
.ends
*
* File: G1_INV1_N2.pex.netlist
* Created: Fri Feb 25 16:24:20 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G1_INV1_N2_VDD 2 5 15 23 28 30 34 37 43 Vss
c22 43 Vss 0.00440656f
c23 34 Vss 7.98732e-19
c24 30 Vss 0.00489873f
c25 28 Vss 0.00252866f
c26 26 Vss 0.00167653f
c27 23 Vss 0.00387287f
c28 15 Vss 0.035607f
c29 14 Vss 0.102409f
c30 5 Vss 0.271444f
r31 34 43 1.16709
r32 32 34 2.41736
r33 31 37 0.326018
r34 30 32 0.652036
r35 30 31 7.46046
r36 26 37 0.326018
r37 26 28 5.50157
r38 23 28 1.16709
r39 17 43 0.0476429
r40 15 17 1.45875
r41 14 18 0.652036
r42 14 17 1.45875
r43 11 15 0.652036
r44 5 18 3.8511
r45 5 11 3.8511
r46 2 23 0.185659
.ends

.subckt PM_G1_INV1_N2_A 2 4 12 22 25 28 Vss
c7 28 Vss 0.00718398f
c8 12 Vss 0.22585f
c9 9 Vss 0.126125f
c10 7 Vss 0.0247918f
c11 4 Vss 0.139046f
r12 22 28 1.16709
r13 22 25 0.0416786
r14 15 28 0.0476429
r15 13 15 0.326018
r16 13 15 0.1167
r17 12 16 0.652036
r18 12 15 6.7686
r19 9 28 0.357321
r20 7 15 0.326018
r21 7 9 0.40845
r22 4 16 3.8511
r23 2 9 3.44265
.ends

.subckt PM_G1_INV1_N2_VSS 3 6 14 24 27 32 37 49 50 56 Vss
c24 51 Vss 0.0012655f
c25 50 Vss 6.56963e-19
c26 49 Vss 0.00353949f
c27 37 Vss 0.00375421f
c28 32 Vss 0.00198022f
c29 27 Vss 2.9624e-19
c30 24 Vss 0.00537236f
c31 15 Vss 0.0358979f
c32 14 Vss 0.0994171f
c33 3 Vss 0.270557f
r34 51 56 0.326018
r35 49 56 0.326018
r36 49 50 7.46046
r37 45 50 0.652036
r38 32 51 5.50157
r39 27 37 1.16709
r40 27 45 2.41736
r41 24 32 1.16709
r42 17 37 0.0476429
r43 15 17 1.45875
r44 14 18 0.652036
r45 14 17 1.45875
r46 11 15 0.652036
r47 6 24 0.185659
r48 3 18 3.8511
r49 3 11 3.8511
.ends

.subckt PM_G1_INV1_N2_Z 2 4 13 16 Vss
c11 13 Vss 0.00523231f
c12 4 Vss 0.00143442f
r13 16 19 0.0416786
r14 13 19 1.16709
r15 4 13 0.185659
r16 2 13 0.185659
.ends

.subckt G1_INV1_N2  VDD A VSS Z
*
* Z	Z
* VSS	VSS
* A	A
* VDD	VDD
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_A_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VDD_XI4.X0_PGD N_A_XI4.X0_CG N_VDD_XI4.X0_PGD
+ N_VSS_XI4.X0_S TIGFET_HPNW8
*
x_PM_G1_INV1_N2_VDD N_VDD_XI6.X0_S N_VDD_XI4.X0_PGD N_VDD_c_4_p N_VDD_c_17_p
+ N_VDD_c_3_p N_VDD_c_5_p N_VDD_c_8_p VDD N_VDD_c_9_p Vss PM_G1_INV1_N2_VDD
x_PM_G1_INV1_N2_A N_A_XI6.X0_CG N_A_XI4.X0_CG N_A_c_23_n N_A_c_25_p A N_A_c_26_p
+ Vss PM_G1_INV1_N2_A
x_PM_G1_INV1_N2_VSS N_VSS_XI6.X0_PGD N_VSS_XI4.X0_S N_VSS_c_32_n N_VSS_c_50_p
+ N_VSS_c_34_n N_VSS_c_38_n N_VSS_c_40_n N_VSS_c_43_n N_VSS_c_44_n VSS Vss
+ PM_G1_INV1_N2_VSS
x_PM_G1_INV1_N2_Z N_Z_XI6.X0_D N_Z_XI4.X0_D N_Z_c_54_n Z Vss PM_G1_INV1_N2_Z
cc_1 N_VDD_XI4.X0_PGD N_A_c_23_n 4.28964e-19
cc_2 N_VDD_XI4.X0_PGD N_VSS_XI6.X0_PGD 0.0020004f
cc_3 N_VDD_c_3_p N_VSS_XI6.X0_PGD 4.31044e-19
cc_4 N_VDD_c_4_p N_VSS_c_32_n 0.0020004f
cc_5 N_VDD_c_5_p N_VSS_c_32_n 5.13652e-19
cc_6 N_VDD_c_3_p N_VSS_c_34_n 0.00287439f
cc_7 N_VDD_c_5_p N_VSS_c_34_n 0.00141709f
cc_8 N_VDD_c_8_p N_VSS_c_34_n 8.61874e-19
cc_9 N_VDD_c_9_p N_VSS_c_34_n 3.48267e-19
cc_10 N_VDD_c_3_p N_VSS_c_38_n 4.56935e-19
cc_11 N_VDD_c_8_p N_VSS_c_38_n 0.00104259f
cc_12 N_VDD_c_3_p N_VSS_c_40_n 9.55109e-19
cc_13 N_VDD_c_5_p N_VSS_c_40_n 0.00103739f
cc_14 N_VDD_c_9_p N_VSS_c_40_n 6.46219e-19
cc_15 N_VDD_c_5_p N_VSS_c_43_n 0.00582834f
cc_16 N_VDD_c_5_p N_VSS_c_44_n 0.00172765f
cc_17 N_VDD_c_17_p N_Z_c_54_n 3.43419e-19
cc_18 N_VDD_c_3_p N_Z_c_54_n 3.48267e-19
cc_19 N_VDD_c_5_p N_Z_c_54_n 3.21105e-19
cc_20 N_VDD_c_17_p Z 3.48267e-19
cc_21 N_VDD_c_3_p Z 7.09569e-19
cc_22 N_VDD_c_5_p Z 4.30066e-19
cc_23 N_A_c_23_n N_VSS_XI6.X0_PGD 4.2599e-19
cc_24 N_A_c_25_p N_VSS_c_34_n 6.08006e-19
cc_25 N_A_c_26_p N_VSS_c_34_n 3.34201e-19
cc_26 N_A_c_25_p N_VSS_c_40_n 3.49905e-19
cc_27 N_A_c_26_p N_VSS_c_40_n 2.68747e-19
cc_28 N_A_c_23_n N_Z_c_54_n 6.55689e-19
cc_29 N_VSS_c_50_p N_Z_c_54_n 3.43419e-19
cc_30 N_VSS_c_38_n N_Z_c_54_n 3.48267e-19
cc_31 N_VSS_c_38_n Z 8.23589e-19
cc_32 N_VSS_c_43_n Z 2.41335e-19
*
.ends
*
*
.subckt INV1_HPNW8 A Y VDD VSS
xgate (VDD A VSS Y) G1_INV1_N2
.ends
*
* File: G3_LATQ1_N2.pex.netlist
* Created: Tue Apr  5 11:38:39 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_LATQ1_N2_VDD 2 4 6 8 10 12 14 16 31 42 44 48 58 63 66 68 69 70 71
+ 72 75 77 81 85 90 92 98 103 Vss
c89 103 Vss 0.00490183f
c90 98 Vss 0.00460926f
c91 90 Vss 2.39889e-19
c92 85 Vss 0.00243594f
c93 83 Vss 0.0016991f
c94 81 Vss 9.06638e-19
c95 77 Vss 0.0042879f
c96 75 Vss 7.26394e-19
c97 72 Vss 8.65068e-19
c98 71 Vss 0.0022063f
c99 70 Vss 8.64091e-19
c100 69 Vss 0.00567616f
c101 68 Vss 0.00905486f
c102 66 Vss 0.00502493f
c103 63 Vss 0.00660615f
c104 58 Vss 0.00394659f
c105 53 Vss 0.0307649f
c106 48 Vss 0.231494f
c107 44 Vss 7.7692e-20
c108 42 Vss 0.0357051f
c109 41 Vss 0.0656875f
c110 32 Vss 0.035919f
c111 31 Vss 0.101295f
c112 16 Vss 0.00143442f
c113 14 Vss 0.137165f
c114 10 Vss 0.136745f
c115 8 Vss 0.135164f
c116 6 Vss 0.13553f
c117 4 Vss 0.135175f
r118 83 92 0.326018
r119 83 85 5.2515
r120 81 103 1.16709
r121 79 81 2.16729
r122 78 90 0.494161
r123 77 92 0.326018
r124 77 78 7.46046
r125 75 98 1.16709
r126 73 90 0.128424
r127 73 75 2.16729
r128 71 90 0.494161
r129 71 72 4.37625
r130 69 79 0.652036
r131 69 70 10.1279
r132 68 72 0.652036
r133 67 68 15.5461
r134 66 89 2.334
r135 66 67 0.14525
r136 65 70 0.652036
r137 65 66 4.62632
r138 63 85 1.16709
r139 58 89 1.16709
r140 49 53 0.494161
r141 48 50 0.652036
r142 48 49 6.8853
r143 45 53 0.128424
r144 44 103 0.0476429
r145 42 44 1.45875
r146 41 53 0.494161
r147 41 44 1.45875
r148 38 42 0.652036
r149 34 98 0.0476429
r150 32 34 1.45875
r151 31 35 0.652036
r152 31 34 1.45875
r153 28 32 0.652036
r154 16 63 0.185659
r155 14 50 3.8511
r156 12 63 0.185659
r157 10 45 3.8511
r158 8 38 3.8511
r159 6 28 3.8511
r160 4 35 3.8511
r161 2 58 0.185659
.ends

.subckt PM_G3_LATQ1_N2_VSS 2 4 6 8 10 12 14 16 31 32 34 42 48 58 63 66 71 76 81
+ 90 95 104 106 107 108 113 114 119 129 130 132 Vss
c81 130 Vss 3.75522e-19
c82 129 Vss 4.28045e-19
c83 125 Vss 0.00128107f
c84 119 Vss 0.00326562f
c85 114 Vss 8.21919e-19
c86 113 Vss 0.00415461f
c87 108 Vss 8.27105e-19
c88 107 Vss 0.00171853f
c89 106 Vss 0.00164009f
c90 104 Vss 0.00508678f
c91 95 Vss 0.00436437f
c92 90 Vss 0.00392783f
c93 81 Vss 0.0023337f
c94 76 Vss 5.9672e-19
c95 71 Vss 4.65089e-19
c96 66 Vss 0.00142325f
c97 63 Vss 0.00655541f
c98 58 Vss 0.00751018f
c99 53 Vss 0.0307649f
c100 48 Vss 0.231624f
c101 42 Vss 0.0348714f
c102 41 Vss 0.0648006f
c103 34 Vss 1.05421e-19
c104 32 Vss 0.0350852f
c105 31 Vss 0.0994129f
c106 16 Vss 0.137353f
c107 14 Vss 0.00143442f
c108 12 Vss 0.137077f
c109 10 Vss 0.135163f
c110 4 Vss 0.135531f
c111 2 Vss 0.135176f
r112 125 132 0.326018
r113 120 130 0.494161
r114 119 132 0.326018
r115 119 120 7.46046
r116 115 130 0.128424
r117 113 121 0.652036
r118 113 114 10.1279
r119 109 129 0.0828784
r120 107 130 0.494161
r121 107 108 4.37625
r122 106 114 0.652036
r123 105 129 0.551426
r124 105 106 4.58464
r125 104 129 0.551426
r126 103 108 0.652036
r127 103 104 15.5878
r128 81 125 5.2515
r129 76 95 1.16709
r130 76 121 2.16729
r131 71 90 1.16709
r132 71 115 2.16729
r133 66 109 1.82344
r134 63 81 1.16709
r135 58 66 1.16709
r136 49 53 0.494161
r137 48 50 0.652036
r138 48 49 6.8853
r139 45 53 0.128424
r140 44 95 0.0476429
r141 42 44 1.45875
r142 41 53 0.494161
r143 41 44 1.45875
r144 38 42 0.652036
r145 34 90 0.0476429
r146 32 34 1.45875
r147 31 35 0.652036
r148 31 34 1.45875
r149 28 32 0.652036
r150 16 50 3.8511
r151 14 63 0.185659
r152 12 45 3.8511
r153 10 38 3.8511
r154 8 63 0.185659
r155 6 58 0.185659
r156 4 28 3.8511
r157 2 35 3.8511
.ends

.subckt PM_G3_LATQ1_N2_G 2 4 6 14 15 22 31 37 Vss
c26 37 Vss 0.00234039f
c27 31 Vss 4.77975e-19
c28 29 Vss 0.0295006f
c29 22 Vss 0.152742f
c30 15 Vss 0.17649f
c31 14 Vss 2.16373e-19
c32 10 Vss 0.0247918f
c33 6 Vss 0.137829f
c34 4 Vss 0.138596f
c35 2 Vss 0.125945f
r36 34 37 1.16709
r37 31 34 0.0833571
r38 23 29 0.494161
r39 22 24 0.652036
r40 22 23 4.84305
r41 19 29 0.128424
r42 18 37 0.0476429
r43 16 18 0.326018
r44 16 18 0.1167
r45 15 29 0.494161
r46 15 18 6.7686
r47 14 37 0.357321
r48 10 18 0.326018
r49 10 14 0.40845
r50 6 24 3.8511
r51 4 19 3.8511
r52 2 14 3.44265
.ends

.subckt PM_G3_LATQ1_N2_QN 2 4 6 8 20 23 33 37 40 45 48 53 69 Vss
c46 69 Vss 4.0109e-19
c47 53 Vss 0.0021144f
c48 48 Vss 0.00823447f
c49 45 Vss 0.00518254f
c50 40 Vss 7.20624e-19
c51 37 Vss 0.00663771f
c52 33 Vss 0.00663771f
c53 23 Vss 2.32346e-19
c54 20 Vss 0.211796f
c55 17 Vss 0.12596f
c56 15 Vss 0.0247918f
c57 4 Vss 0.137276f
r58 65 69 0.652036
r59 48 69 13.7956
r60 48 50 5.50157
r61 45 48 5.50157
r62 40 53 1.16709
r63 40 65 1.83386
r64 37 50 1.16709
r65 33 45 1.16709
r66 23 53 0.0476429
r67 21 23 0.326018
r68 21 23 0.1167
r69 20 24 0.652036
r70 20 23 6.7686
r71 17 53 0.357321
r72 15 23 0.326018
r73 15 17 0.40845
r74 8 37 0.185659
r75 6 33 0.185659
r76 4 24 3.8511
r77 2 17 3.44265
.ends

.subckt PM_G3_LATQ1_N2_GN 2 4 6 12 23 27 29 30 32 39 Vss
c44 39 Vss 0.0045172f
c45 32 Vss 8.57161e-19
c46 30 Vss 7.68504e-19
c47 29 Vss 0.00117249f
c48 27 Vss 0.00109299f
c49 23 Vss 0.00551775f
c50 12 Vss 0.171663f
c51 6 Vss 0.232172f
c52 4 Vss 0.00143442f
r53 32 39 1.16709
r54 29 32 0.531835
r55 29 30 1.70882
r56 25 30 0.652036
r57 25 27 4.91807
r58 23 27 1.16709
r59 14 39 0.197068
r60 12 16 0.652036
r61 12 14 4.668
r62 6 16 7.1187
r63 4 23 0.185659
r64 2 23 0.185659
.ends

.subckt PM_G3_LATQ1_N2_Q 2 4 13 18 Vss
c12 18 Vss 3.58669e-19
c13 13 Vss 0.004507f
c14 4 Vss 0.00143442f
r15 13 18 1.16709
r16 4 13 0.185659
r17 2 13 0.185659
.ends

.subckt PM_G3_LATQ1_N2_D 2 4 10 14 Vss
c14 14 Vss 4.15825e-19
c15 10 Vss 1.35847e-19
c16 2 Vss 0.475046f
r17 14 17 0.0416786
r18 10 17 1.16709
r19 4 10 7.7022
r20 2 10 7.7022
.ends

.subckt G3_LATQ1_N2  VDD VSS G Q D
*
* D	D
* Q	Q
* G	G
* VSS	VSS
* VDD	VDD
XI6.X0 N_GN_XI6.X0_D N_VSS_XI6.X0_PGD N_G_XI6.X0_CG N_VSS_XI6.X0_PGS
+ N_VDD_XI6.X0_S TIGFET_HPNW8
XI10.X0 N_Q_XI10.X0_D N_VDD_XI10.X0_PGD N_QN_XI10.X0_CG N_VDD_XI10.X0_PGS
+ N_VSS_XI10.X0_S TIGFET_HPNW8
XI9.X0 N_GN_XI9.X0_D N_VDD_XI9.X0_PGD N_G_XI9.X0_CG N_VDD_XI9.X0_PGS
+ N_VSS_XI9.X0_S TIGFET_HPNW8
XI8.X0 N_Q_XI8.X0_D N_VSS_XI8.X0_PGD N_QN_XI8.X0_CG N_VSS_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW8
XI11.X0 N_QN_XI11.X0_D N_VDD_XI11.X0_PGD N_D_XI11.X0_CG N_G_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW8
XI7.X0 N_QN_XI7.X0_D N_VSS_XI7.X0_PGD N_D_XI7.X0_CG N_GN_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW8
*
x_PM_G3_LATQ1_N2_VDD N_VDD_XI6.X0_S N_VDD_XI10.X0_PGD N_VDD_XI10.X0_PGS
+ N_VDD_XI9.X0_PGD N_VDD_XI9.X0_PGS N_VDD_XI8.X0_S N_VDD_XI11.X0_PGD
+ N_VDD_XI7.X0_S N_VDD_c_9_p N_VDD_c_5_p N_VDD_c_81_p N_VDD_c_15_p N_VDD_c_13_p
+ N_VDD_c_11_p N_VDD_c_7_p N_VDD_c_14_p N_VDD_c_6_p N_VDD_c_42_p N_VDD_c_19_p
+ N_VDD_c_46_p N_VDD_c_24_p N_VDD_c_10_p N_VDD_c_22_p N_VDD_c_12_p N_VDD_c_45_p
+ VDD N_VDD_c_27_p N_VDD_c_23_p Vss PM_G3_LATQ1_N2_VDD
x_PM_G3_LATQ1_N2_VSS N_VSS_XI6.X0_PGD N_VSS_XI6.X0_PGS N_VSS_XI10.X0_S
+ N_VSS_XI9.X0_S N_VSS_XI8.X0_PGD N_VSS_XI8.X0_PGS N_VSS_XI11.X0_S
+ N_VSS_XI7.X0_PGD N_VSS_c_94_n N_VSS_c_96_n N_VSS_c_139_p N_VSS_c_98_n
+ N_VSS_c_100_n N_VSS_c_102_n N_VSS_c_104_n N_VSS_c_106_n N_VSS_c_109_n
+ N_VSS_c_113_n N_VSS_c_117_n N_VSS_c_119_n N_VSS_c_123_n N_VSS_c_127_n
+ N_VSS_c_129_n N_VSS_c_130_n N_VSS_c_131_n N_VSS_c_132_n N_VSS_c_135_n
+ N_VSS_c_136_n N_VSS_c_137_n N_VSS_c_138_n VSS Vss PM_G3_LATQ1_N2_VSS
x_PM_G3_LATQ1_N2_G N_G_XI6.X0_CG N_G_XI9.X0_CG N_G_XI11.X0_PGS N_G_c_176_n
+ N_G_c_172_n N_G_c_173_n G N_G_c_175_n Vss PM_G3_LATQ1_N2_G
x_PM_G3_LATQ1_N2_QN N_QN_XI10.X0_CG N_QN_XI8.X0_CG N_QN_XI11.X0_D N_QN_XI7.X0_D
+ N_QN_c_197_n N_QN_c_198_n N_QN_c_214_n N_QN_c_199_n N_QN_c_201_n N_QN_c_204_n
+ N_QN_c_206_n N_QN_c_209_n N_QN_c_212_n Vss PM_G3_LATQ1_N2_QN
x_PM_G3_LATQ1_N2_GN N_GN_XI6.X0_D N_GN_XI9.X0_D N_GN_XI7.X0_PGS N_GN_c_243_n
+ N_GN_c_246_n N_GN_c_249_n N_GN_c_269_n N_GN_c_275_n N_GN_c_276_n N_GN_c_253_n
+ Vss PM_G3_LATQ1_N2_GN
x_PM_G3_LATQ1_N2_Q N_Q_XI10.X0_D N_Q_XI8.X0_D N_Q_c_287_n Q Vss PM_G3_LATQ1_N2_Q
x_PM_G3_LATQ1_N2_D N_D_XI11.X0_CG N_D_XI7.X0_CG N_D_c_304_n D Vss
+ PM_G3_LATQ1_N2_D
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI6.X0_PGD 0.00203852f
cc_2 N_VDD_XI10.X0_PGS N_VSS_XI6.X0_PGS 2.37403e-19
cc_3 N_VDD_XI10.X0_PGD N_VSS_XI8.X0_PGD 0.00203076f
cc_4 N_VDD_XI11.X0_PGD N_VSS_XI7.X0_PGD 2.37403e-19
cc_5 N_VDD_c_5_p N_VSS_c_94_n 0.00203852f
cc_6 N_VDD_c_6_p N_VSS_c_94_n 3.9313e-19
cc_7 N_VDD_c_7_p N_VSS_c_96_n 3.80615e-19
cc_8 N_VDD_c_6_p N_VSS_c_96_n 3.9313e-19
cc_9 N_VDD_c_9_p N_VSS_c_98_n 0.00203076f
cc_10 N_VDD_c_10_p N_VSS_c_98_n 2.95583e-19
cc_11 N_VDD_c_11_p N_VSS_c_100_n 2.64155e-19
cc_12 N_VDD_c_12_p N_VSS_c_100_n 8.58125e-19
cc_13 N_VDD_c_13_p N_VSS_c_102_n 2.12761e-19
cc_14 N_VDD_c_14_p N_VSS_c_102_n 9.5668e-19
cc_15 N_VDD_c_15_p N_VSS_c_104_n 2.64155e-19
cc_16 N_VDD_c_11_p N_VSS_c_104_n 2.69828e-19
cc_17 N_VDD_c_7_p N_VSS_c_106_n 4.61436e-19
cc_18 N_VDD_c_14_p N_VSS_c_106_n 0.00165395f
cc_19 N_VDD_c_19_p N_VSS_c_106_n 4.5625e-19
cc_20 N_VDD_c_7_p N_VSS_c_109_n 9.31121e-19
cc_21 N_VDD_c_6_p N_VSS_c_109_n 0.00161703f
cc_22 N_VDD_c_22_p N_VSS_c_109_n 7.09654e-19
cc_23 N_VDD_c_23_p N_VSS_c_109_n 3.48267e-19
cc_24 N_VDD_c_24_p N_VSS_c_113_n 9.52068e-19
cc_25 N_VDD_c_10_p N_VSS_c_113_n 0.00141228f
cc_26 N_VDD_c_12_p N_VSS_c_113_n 0.00257912f
cc_27 N_VDD_c_27_p N_VSS_c_113_n 3.48267e-19
cc_28 N_VDD_c_7_p N_VSS_c_117_n 2.12713e-19
cc_29 N_VDD_c_22_p N_VSS_c_117_n 8.43845e-19
cc_30 N_VDD_c_7_p N_VSS_c_119_n 4.24454e-19
cc_31 N_VDD_c_6_p N_VSS_c_119_n 2.26455e-19
cc_32 N_VDD_c_22_p N_VSS_c_119_n 3.84769e-19
cc_33 N_VDD_c_23_p N_VSS_c_119_n 6.489e-19
cc_34 N_VDD_c_24_p N_VSS_c_123_n 3.82294e-19
cc_35 N_VDD_c_10_p N_VSS_c_123_n 0.00114511f
cc_36 N_VDD_c_12_p N_VSS_c_123_n 9.55109e-19
cc_37 N_VDD_c_27_p N_VSS_c_123_n 6.46219e-19
cc_38 N_VDD_c_7_p N_VSS_c_127_n 0.00468852f
cc_39 N_VDD_c_14_p N_VSS_c_127_n 0.00657271f
cc_40 N_VDD_c_14_p N_VSS_c_129_n 0.00377187f
cc_41 N_VDD_c_6_p N_VSS_c_130_n 0.00345737f
cc_42 N_VDD_c_42_p N_VSS_c_131_n 0.00106538f
cc_43 N_VDD_c_19_p N_VSS_c_132_n 0.00353938f
cc_44 N_VDD_c_10_p N_VSS_c_132_n 0.00581493f
cc_45 N_VDD_c_45_p N_VSS_c_132_n 9.99051e-19
cc_46 N_VDD_c_46_p N_VSS_c_135_n 0.0010616f
cc_47 N_VDD_c_6_p N_VSS_c_136_n 0.00566938f
cc_48 N_VDD_c_14_p N_VSS_c_137_n 9.16632e-19
cc_49 N_VDD_c_6_p N_VSS_c_138_n 7.74609e-19
cc_50 N_VDD_c_15_p N_G_XI11.X0_PGS 0.00163289f
cc_51 N_VDD_XI9.X0_PGD N_G_c_172_n 3.96934e-19
cc_52 N_VDD_XI9.X0_PGS N_G_c_173_n 4.08222e-19
cc_53 N_VDD_c_14_p G 5.04211e-19
cc_54 N_VDD_c_14_p N_G_c_175_n 5.56409e-19
cc_55 N_VDD_XI10.X0_PGD N_QN_c_197_n 4.07423e-19
cc_56 N_VDD_c_27_p N_QN_c_198_n 0.00100159f
cc_57 N_VDD_c_11_p N_QN_c_199_n 3.43419e-19
cc_58 N_VDD_c_12_p N_QN_c_199_n 3.48267e-19
cc_59 N_VDD_c_14_p N_QN_c_201_n 4.08289e-19
cc_60 N_VDD_c_24_p N_QN_c_201_n 2.98644e-19
cc_61 N_VDD_c_27_p N_QN_c_201_n 3.15998e-19
cc_62 N_VDD_c_11_p N_QN_c_204_n 3.48267e-19
cc_63 N_VDD_c_12_p N_QN_c_204_n 9.04108e-19
cc_64 N_VDD_c_6_p N_QN_c_206_n 3.90695e-19
cc_65 N_VDD_c_10_p N_QN_c_206_n 3.49463e-19
cc_66 N_VDD_c_12_p N_QN_c_206_n 3.67848e-19
cc_67 N_VDD_c_14_p N_QN_c_209_n 6.60137e-19
cc_68 N_VDD_c_24_p N_QN_c_209_n 3.43988e-19
cc_69 N_VDD_c_27_p N_QN_c_209_n 2.68747e-19
cc_70 N_VDD_c_14_p N_QN_c_212_n 3.90734e-19
cc_71 N_VDD_XI9.X0_PGS N_GN_c_243_n 3.40745e-19
cc_72 N_VDD_c_15_p N_GN_c_243_n 2.49684e-19
cc_73 N_VDD_c_11_p N_GN_c_243_n 3.08361e-19
cc_74 N_VDD_c_13_p N_GN_c_246_n 3.43419e-19
cc_75 N_VDD_c_7_p N_GN_c_246_n 3.72199e-19
cc_76 N_VDD_c_6_p N_GN_c_246_n 3.4118e-19
cc_77 N_VDD_c_13_p N_GN_c_249_n 3.48267e-19
cc_78 N_VDD_c_7_p N_GN_c_249_n 7.94301e-19
cc_79 N_VDD_c_14_p N_GN_c_249_n 0.0010243f
cc_80 N_VDD_c_6_p N_GN_c_249_n 4.77682e-19
cc_81 N_VDD_c_81_p N_GN_c_253_n 3.88849e-19
cc_82 N_VDD_c_22_p N_GN_c_253_n 2.02851e-19
cc_83 N_VDD_c_11_p N_Q_c_287_n 3.43419e-19
cc_84 N_VDD_c_10_p N_Q_c_287_n 3.4118e-19
cc_85 N_VDD_c_12_p N_Q_c_287_n 3.48267e-19
cc_86 N_VDD_c_11_p Q 3.48267e-19
cc_87 N_VDD_c_10_p Q 4.58391e-19
cc_88 N_VDD_c_12_p Q 7.09569e-19
cc_89 N_VDD_c_15_p N_D_XI11.X0_CG 4.20341e-19
cc_90 N_VSS_c_139_p N_G_c_176_n 9.37683e-19
cc_91 N_VSS_XI6.X0_PGD N_G_c_172_n 4.04227e-19
cc_92 N_VSS_c_109_n G 3.00355e-19
cc_93 N_VSS_c_119_n G 3.2351e-19
cc_94 N_VSS_c_127_n G 2.86445e-19
cc_95 N_VSS_c_109_n N_G_c_175_n 3.2351e-19
cc_96 N_VSS_c_119_n N_G_c_175_n 2.68747e-19
cc_97 N_VSS_XI8.X0_PGD N_QN_c_197_n 3.93738e-19
cc_98 N_VSS_c_104_n N_QN_c_214_n 3.43419e-19
cc_99 N_VSS_c_117_n N_QN_c_214_n 3.48267e-19
cc_100 N_VSS_c_132_n N_QN_c_201_n 2.32769e-19
cc_101 N_VSS_c_104_n N_QN_c_204_n 3.48267e-19
cc_102 N_VSS_c_117_n N_QN_c_204_n 8.62542e-19
cc_103 N_VSS_c_113_n N_QN_c_206_n 2.72578e-19
cc_104 N_VSS_c_117_n N_QN_c_206_n 6.59201e-19
cc_105 N_VSS_c_132_n N_QN_c_206_n 5.73383e-19
cc_106 N_VSS_c_136_n N_QN_c_206_n 7.86339e-19
cc_107 N_VSS_c_109_n N_QN_c_212_n 4.50267e-19
cc_108 N_VSS_c_127_n N_QN_c_212_n 0.00182171f
cc_109 N_VSS_c_100_n N_GN_XI7.X0_PGS 0.00172633f
cc_110 N_VSS_XI8.X0_PGS N_GN_c_243_n 6.82193e-19
cc_111 N_VSS_c_104_n N_GN_c_246_n 3.43419e-19
cc_112 N_VSS_c_117_n N_GN_c_246_n 3.48267e-19
cc_113 N_VSS_c_104_n N_GN_c_249_n 3.48267e-19
cc_114 N_VSS_c_117_n N_GN_c_249_n 4.99861e-19
cc_115 N_VSS_c_127_n N_GN_c_249_n 5.59824e-19
cc_116 N_VSS_c_113_n N_GN_c_253_n 2.02167e-19
cc_117 N_VSS_c_123_n N_GN_c_253_n 3.56129e-19
cc_118 N_VSS_c_102_n N_Q_c_287_n 3.43419e-19
cc_119 N_VSS_c_106_n N_Q_c_287_n 3.48267e-19
cc_120 N_VSS_c_106_n Q 8.15956e-19
cc_121 N_VSS_c_100_n N_D_XI11.X0_CG 4.20341e-19
cc_122 N_G_c_172_n N_QN_c_197_n 0.00398811f
cc_123 G N_QN_c_201_n 4.48861e-19
cc_124 N_G_c_175_n N_QN_c_201_n 4.54925e-19
cc_125 G N_QN_c_209_n 4.56568e-19
cc_126 N_G_c_175_n N_QN_c_209_n 0.00268575f
cc_127 N_G_c_173_n N_GN_c_243_n 0.00842907f
cc_128 N_G_c_172_n N_GN_c_246_n 6.8653e-19
cc_129 N_G_c_172_n N_GN_c_249_n 3.82175e-19
cc_130 G N_GN_c_249_n 0.00151253f
cc_131 N_G_c_175_n N_GN_c_249_n 9.72448e-19
cc_132 N_G_c_172_n N_GN_c_269_n 3.75306e-19
cc_133 N_G_c_172_n N_GN_c_253_n 0.00395135f
cc_134 N_G_c_175_n N_GN_c_253_n 2.41671e-19
cc_135 N_G_XI11.X0_PGS N_D_XI11.X0_CG 0.00435077f
cc_136 N_QN_c_197_n N_GN_XI7.X0_PGS 0.00196434f
cc_137 N_QN_c_204_n N_GN_c_249_n 0.0010213f
cc_138 N_QN_c_206_n N_GN_c_269_n 9.45997e-19
cc_139 N_QN_c_206_n N_GN_c_275_n 0.00125885f
cc_140 N_QN_c_206_n N_GN_c_276_n 9.71021e-19
cc_141 N_QN_c_197_n N_GN_c_253_n 0.00340055f
cc_142 N_QN_c_209_n N_GN_c_253_n 2.75519e-19
cc_143 N_QN_c_197_n N_Q_c_287_n 6.8653e-19
cc_144 N_QN_c_197_n N_D_XI11.X0_CG 3.26559e-19
cc_145 N_QN_c_204_n N_D_XI11.X0_CG 0.0010503f
cc_146 N_QN_c_204_n N_D_c_304_n 0.00130556f
cc_147 N_QN_c_204_n D 0.00141415f
cc_148 N_QN_c_206_n D 0.00146947f
cc_149 N_GN_c_275_n N_Q_c_287_n 4.09054e-19
cc_150 N_GN_c_275_n Q 5.11868e-19
cc_151 N_GN_XI7.X0_PGS N_D_XI11.X0_CG 0.0048787f
cc_152 N_GN_c_243_n N_D_c_304_n 0.00333193f
cc_153 N_GN_c_276_n N_D_c_304_n 3.73302e-19
cc_154 N_GN_c_253_n N_D_c_304_n 8.5422e-19
cc_155 N_GN_c_276_n D 2.85187e-19
cc_156 N_GN_c_253_n D 3.48267e-19
*
.ends
*
*
.subckt LATQ1_HPNW8 D G Q VDD VSS
xgate (VDD VSS G Q D) G3_LATQ1_N2
.ends
*
* File: G4_MAJ3_N2.pex.netlist
* Created: Fri Mar  4 11:26:54 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MAJ3_N2_VDD 2 4 7 11 27 28 30 31 32 44 48 52 54 56 57 58 61 63 67
+ 69 70 73 77 79 80 90 95 Vss
c77 95 Vss 0.00486523f
c78 90 Vss 0.00461066f
c79 80 Vss 4.52364e-19
c80 79 Vss 4.28405e-19
c81 77 Vss 4.66438e-19
c82 73 Vss 8.57616e-19
c83 70 Vss 8.64091e-19
c84 69 Vss 0.00558016f
c85 67 Vss 0.00139758f
c86 63 Vss 0.00140124f
c87 58 Vss 8.64091e-19
c88 57 Vss 0.00559492f
c89 56 Vss 0.00209681f
c90 54 Vss 0.00571364f
c91 52 Vss 0.00207954f
c92 48 Vss 0.00382489f
c93 44 Vss 0.00532438f
c94 32 Vss 0.035607f
c95 31 Vss 0.100823f
c96 28 Vss 0.035607f
c97 27 Vss 0.100961f
c98 11 Vss 0.266772f
c99 7 Vss 0.268336f
r100 77 95 1.16709
r101 75 77 2.16729
r102 73 90 1.16709
r103 71 73 2.16729
r104 69 75 0.652036
r105 69 70 10.1279
r106 65 80 0.0828784
r107 65 67 1.82344
r108 61 63 1.167
r109 59 79 0.0828784
r110 59 61 0.656438
r111 57 71 0.652036
r112 57 58 10.1279
r113 56 70 0.652036
r114 55 80 0.551426
r115 55 56 4.58464
r116 54 80 0.551426
r117 53 79 0.551426
r118 53 54 9.66943
r119 52 79 0.551426
r120 51 58 0.652036
r121 51 52 4.58464
r122 48 67 1.16709
r123 44 63 1.16709
r124 34 95 0.0476429
r125 32 34 1.45875
r126 31 38 0.652036
r127 31 34 1.45875
r128 30 90 0.0476429
r129 28 30 1.45875
r130 27 35 0.652036
r131 27 30 1.45875
r132 24 32 0.652036
r133 21 28 0.652036
r134 11 38 3.8511
r135 11 24 3.8511
r136 7 35 3.8511
r137 7 21 3.8511
r138 4 48 0.185659
r139 2 44 0.185659
.ends

.subckt PM_G4_MAJ3_N2_VSS 3 7 10 12 27 28 30 31 32 45 49 52 57 62 67 70 73 78 91
+ 92 93 94 95 104 114 115 117 Vss
c83 115 Vss 3.75522e-19
c84 114 Vss 3.75522e-19
c85 110 Vss 0.00128107f
c86 104 Vss 0.00335813f
c87 95 Vss 8.27105e-19
c88 94 Vss 0.00156442f
c89 93 Vss 8.27105e-19
c90 92 Vss 0.00156442f
c91 91 Vss 0.00686995f
c92 78 Vss 0.00393332f
c93 73 Vss 0.00431768f
c94 70 Vss 0.00351391f
c95 67 Vss 0.00277973f
c96 62 Vss 0.00186148f
c97 57 Vss 0.00131291f
c98 52 Vss 0.00112626f
c99 49 Vss 0.00527641f
c100 45 Vss 0.00377692f
c101 32 Vss 0.0350852f
c102 31 Vss 0.0994129f
c103 30 Vss 9.50876e-20
c104 28 Vss 0.0350852f
c105 27 Vss 0.0994129f
c106 7 Vss 0.267138f
c107 3 Vss 0.268863f
r108 110 117 0.326018
r109 106 115 0.494161
r110 105 114 0.494161
r111 104 117 0.326018
r112 104 105 7.46046
r113 100 115 0.128424
r114 96 114 0.128424
r115 94 115 0.494161
r116 94 95 4.37625
r117 92 114 0.494161
r118 92 93 4.37625
r119 91 95 0.652036
r120 90 93 0.652036
r121 90 91 21.5061
r122 70 106 8.04396
r123 67 70 5.835
r124 62 110 5.2515
r125 57 78 1.16709
r126 57 100 2.16729
r127 52 73 1.16709
r128 52 96 2.16729
r129 49 67 1.16709
r130 45 62 1.16709
r131 34 78 0.0476429
r132 32 34 1.45875
r133 31 38 0.652036
r134 31 34 1.45875
r135 30 73 0.0476429
r136 28 30 1.45875
r137 27 35 0.652036
r138 27 30 1.45875
r139 24 32 0.652036
r140 21 28 0.652036
r141 12 49 0.185659
r142 10 45 0.185659
r143 7 38 3.8511
r144 7 24 3.8511
r145 3 35 3.8511
r146 3 21 3.8511
.ends

.subckt PM_G4_MAJ3_N2_A 1 2 4 6 9 13 31 53 57 62 67 71 74 76 78 81 89 91 99 100
+ 102 111 Vss
c78 111 Vss 0.00528881f
c79 102 Vss 0.00500597f
c80 99 Vss 0.00422425f
c81 96 Vss 7.53731e-19
c82 91 Vss 7.84512e-19
c83 89 Vss 8.92851e-19
c84 85 Vss 0.00253152f
c85 81 Vss 7.20282e-19
c86 78 Vss 0.0011176f
c87 77 Vss 0.00146569f
c88 76 Vss 0.00441934f
c89 71 Vss 0.00722904f
c90 67 Vss 0.00399277f
c91 62 Vss 0.00496845f
c92 57 Vss 0.135055f
c93 53 Vss 0.12803f
c94 31 Vss 0.215113f
c95 27 Vss 0.126125f
c96 25 Vss 0.0247918f
c97 9 Vss 1.22732f
c98 2 Vss 0.139046f
r99 111 114 0.1
r100 98 111 1.16709
r101 98 100 0.490235
r102 98 99 0.490235
r103 94 102 1.16709
r104 91 94 1.08364
r105 87 89 2.50071
r106 85 87 0.653045
r107 85 100 1.5949
r108 84 96 0.466409
r109 84 99 6.9631
r110 79 96 0.152298
r111 79 81 2.50071
r112 77 96 0.466409
r113 77 78 1.7116
r114 75 78 0.653045
r115 75 76 8.7525
r116 72 91 0.0685365
r117 72 74 1.45875
r118 71 76 0.652036
r119 71 74 8.7525
r120 67 89 1.16709
r121 62 81 1.16709
r122 55 57 4.53833
r123 52 114 0.0238214
r124 52 53 2.26917
r125 49 52 2.26917
r126 44 57 0.00605528
r127 43 53 0.00605528
r128 40 55 0.00605528
r129 39 49 0.00605528
r130 34 102 0.0476429
r131 32 34 0.326018
r132 32 34 0.1167
r133 31 35 0.652036
r134 31 34 6.7686
r135 27 102 0.357321
r136 25 34 0.326018
r137 25 27 0.40845
r138 13 44 3.8511
r139 13 40 3.8511
r140 9 13 15.4044
r141 9 43 3.8511
r142 9 13 15.4044
r143 9 39 3.8511
r144 6 67 0.185659
r145 4 62 0.185659
r146 2 35 3.8511
r147 1 27 3.44265
.ends

.subckt PM_G4_MAJ3_N2_BI 2 4 5 6 20 29 34 39 44 54 59 68 74 75 83 Vss
c58 83 Vss 4.27892e-19
c59 75 Vss 3.15444e-19
c60 74 Vss 7.27663e-19
c61 68 Vss 0.00155105f
c62 59 Vss 0.00147096f
c63 54 Vss 0.00139826f
c64 44 Vss 0.00152385f
c65 39 Vss 0.00577944f
c66 34 Vss 0.00175738f
c67 29 Vss 0.00439389f
c68 20 Vss 0.111942f
c69 5 Vss 0.111942f
c70 4 Vss 0.00143442f
r71 79 83 0.655813
r72 74 75 0.65228
r73 73 74 3.42052
r74 68 73 0.65409
r75 44 59 1.16709
r76 44 75 2.1395
r77 39 54 1.16709
r78 39 83 12.0712
r79 39 68 1.96931
r80 34 51 1.16709
r81 34 79 2.334
r82 29 51 0.1
r83 20 59 0.50025
r84 17 54 0.50025
r85 6 20 3.09255
r86 5 17 3.09255
r87 4 29 0.185659
r88 2 29 0.185659
.ends

.subckt PM_G4_MAJ3_N2_AI 2 4 7 11 31 37 43 46 51 60 69 Vss
c44 69 Vss 4.10597e-19
c45 60 Vss 0.00527726f
c46 51 Vss 0.00584502f
c47 46 Vss 0.00110084f
c48 43 Vss 0.00447686f
c49 37 Vss 0.127877f
c50 31 Vss 0.134503f
c51 7 Vss 1.21876f
c52 4 Vss 0.00143442f
r53 65 69 0.652036
r54 60 63 0.1
r55 51 63 1.16709
r56 51 69 13.7539
r57 46 65 2.58407
r58 43 46 1.16709
r59 36 60 0.0238214
r60 36 37 2.334
r61 33 36 2.20433
r62 29 31 4.53833
r63 26 37 0.00605528
r64 25 31 0.00605528
r65 22 33 0.00605528
r66 21 29 0.00605528
r67 11 26 3.8511
r68 11 22 3.8511
r69 7 11 15.4044
r70 7 25 3.8511
r71 7 11 15.4044
r72 7 21 3.8511
r73 4 43 0.185659
r74 2 43 0.185659
.ends

.subckt PM_G4_MAJ3_N2_B 1 2 3 4 13 14 24 42 46 49 54 59 64 69 77 78 84 91 96 97
+ Vss
c68 97 Vss 4.67818e-19
c69 96 Vss 0.00212566f
c70 91 Vss 9.32419e-19
c71 84 Vss 5.17496e-19
c72 78 Vss 3.17701e-19
c73 77 Vss 0.00357974f
c74 69 Vss 0.00148026f
c75 64 Vss 0.0010348f
c76 59 Vss 0.00464385f
c77 54 Vss 0.00163559f
c78 49 Vss 7.01001e-19
c79 46 Vss 5.25457e-19
c80 42 Vss 5.46753e-19
c81 24 Vss 0.111942f
c82 17 Vss 0.0247918f
c83 14 Vss 0.0349292f
c84 13 Vss 0.183407f
c85 4 Vss 0.111942f
c86 2 Vss 0.111095f
c87 1 Vss 0.118069f
r88 95 97 0.65409
r89 95 96 3.42052
r90 91 96 0.65228
r91 87 91 2.1006
r92 84 87 2.04225
r93 77 84 0.0685365
r94 77 78 10.3363
r95 73 78 0.652036
r96 54 69 1.16709
r97 54 97 2.00578
r98 49 64 1.16709
r99 49 87 0.0416786
r100 42 59 1.16709
r101 42 73 2.16729
r102 42 46 0.0530455
r103 36 59 0.238214
r104 33 69 0.50025
r105 24 64 0.50025
r106 22 36 0.262036
r107 17 36 0.326018
r108 17 22 0.05835
r109 14 36 6.7686
r110 13 36 0.326018
r111 13 36 0.1167
r112 9 14 0.652036
r113 4 33 3.09255
r114 3 24 3.09255
r115 2 22 3.09255
r116 1 9 3.1509
.ends

.subckt PM_G4_MAJ3_N2_C 2 4 12 17 20 25 51 Vss
c18 25 Vss 0.00550018f
c19 20 Vss 7.32915e-19
c20 17 Vss 0.00502472f
c21 12 Vss 0.00387713f
r22 25 51 1.78697
r23 20 51 8.27841
r24 17 25 1.16709
r25 12 20 1.16709
r26 4 17 0.185659
r27 2 12 0.185659
.ends

.subckt PM_G4_MAJ3_N2_Z 2 4 6 8 23 27 30 33 Vss
c30 30 Vss 0.00298505f
c31 27 Vss 0.00857889f
c32 23 Vss 0.00745393f
c33 8 Vss 0.00143442f
c34 6 Vss 0.00143442f
r35 33 35 6.04339
r36 30 33 4.95975
r37 27 35 1.16709
r38 23 30 1.16709
r39 8 27 0.185659
r40 6 23 0.185659
r41 4 27 0.185659
r42 2 23 0.185659
.ends

.subckt G4_MAJ3_N2  VDD VSS A B C Z
*
* Z	Z
* C	C
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI11.X0 N_BI_XI11.X0_D N_VSS_XI11.X0_PGD N_B_XI11.X0_CG N_VSS_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW8
XI10.X0 N_AI_XI10.X0_D N_VSS_XI10.X0_PGD N_A_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW8
XI9.X0 N_BI_XI9.X0_D N_VDD_XI9.X0_PGD N_B_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW8
XI0.X0 N_AI_XI0.X0_D N_VDD_XI0.X0_PGD N_A_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_AI_XI15.X0_PGD N_BI_XI15.X0_CG N_AI_XI15.X0_PGD
+ N_A_XI15.X0_S TIGFET_HPNW8
XI13.X0 N_Z_XI13.X0_D N_AI_XI13.X0_PGD N_B_XI13.X0_CG N_AI_XI13.X0_PGD
+ N_C_XI13.X0_S TIGFET_HPNW8
XI14.X0 N_Z_XI14.X0_D N_A_XI14.X0_PGD N_B_XI14.X0_CG N_A_XI14.X0_PGD
+ N_A_XI14.X0_S TIGFET_HPNW8
XI12.X0 N_Z_XI12.X0_D N_A_XI12.X0_PGD N_BI_XI12.X0_CG N_A_XI12.X0_PGD
+ N_C_XI12.X0_S TIGFET_HPNW8
*
x_PM_G4_MAJ3_N2_VDD N_VDD_XI11.X0_S N_VDD_XI10.X0_S N_VDD_XI9.X0_PGD
+ N_VDD_XI0.X0_PGD N_VDD_c_62_p N_VDD_c_4_p N_VDD_c_72_p N_VDD_c_63_p
+ N_VDD_c_8_p N_VDD_c_55_p N_VDD_c_64_p N_VDD_c_6_p N_VDD_c_32_p N_VDD_c_3_p
+ N_VDD_c_5_p N_VDD_c_38_p VDD N_VDD_c_37_p N_VDD_c_39_p N_VDD_c_9_p
+ N_VDD_c_41_p N_VDD_c_13_p N_VDD_c_17_p N_VDD_c_34_p N_VDD_c_35_p N_VDD_c_14_p
+ N_VDD_c_18_p Vss PM_G4_MAJ3_N2_VDD
x_PM_G4_MAJ3_N2_VSS N_VSS_XI11.X0_PGD N_VSS_XI10.X0_PGD N_VSS_XI9.X0_S
+ N_VSS_XI0.X0_S N_VSS_c_81_n N_VSS_c_83_n N_VSS_c_135_p N_VSS_c_85_n
+ N_VSS_c_87_n N_VSS_c_123_p N_VSS_c_125_p N_VSS_c_88_n N_VSS_c_92_n
+ N_VSS_c_96_n N_VSS_c_97_n N_VSS_c_100_n N_VSS_c_101_n N_VSS_c_105_n
+ N_VSS_c_108_n N_VSS_c_113_n N_VSS_c_115_n N_VSS_c_116_n N_VSS_c_118_n
+ N_VSS_c_119_n N_VSS_c_120_n N_VSS_c_121_n VSS Vss PM_G4_MAJ3_N2_VSS
x_PM_G4_MAJ3_N2_A N_A_XI10.X0_CG N_A_XI0.X0_CG N_A_XI15.X0_S N_A_XI14.X0_S
+ N_A_XI14.X0_PGD N_A_XI12.X0_PGD N_A_c_161_n N_A_c_201_p N_A_c_203_p
+ N_A_c_172_n N_A_c_228_p N_A_c_162_n A N_A_c_179_n N_A_c_167_n N_A_c_223_p
+ N_A_c_230_p N_A_c_169_n N_A_c_187_p N_A_c_215_p N_A_c_170_n N_A_c_216_p Vss
+ PM_G4_MAJ3_N2_A
x_PM_G4_MAJ3_N2_BI N_BI_XI11.X0_D N_BI_XI9.X0_D N_BI_XI15.X0_CG N_BI_XI12.X0_CG
+ N_BI_c_252_n N_BI_c_239_n N_BI_c_241_n N_BI_c_249_n N_BI_c_257_n N_BI_c_258_n
+ N_BI_c_259_n N_BI_c_260_n N_BI_c_280_p N_BI_c_283_p N_BI_c_261_n Vss
+ PM_G4_MAJ3_N2_BI
x_PM_G4_MAJ3_N2_AI N_AI_XI10.X0_D N_AI_XI0.X0_D N_AI_XI15.X0_PGD
+ N_AI_XI13.X0_PGD N_AI_c_299_n N_AI_c_300_n N_AI_c_301_n N_AI_c_303_n
+ N_AI_c_306_n N_AI_c_315_n N_AI_c_316_n Vss PM_G4_MAJ3_N2_AI
x_PM_G4_MAJ3_N2_B N_B_XI11.X0_CG N_B_XI9.X0_CG N_B_XI13.X0_CG N_B_XI14.X0_CG
+ N_B_c_341_n N_B_c_355_n N_B_c_393_n N_B_c_342_n B N_B_c_374_n N_B_c_359_n
+ N_B_c_346_n N_B_c_378_n N_B_c_364_n N_B_c_351_n N_B_c_370_n N_B_c_371_n
+ N_B_c_387_n N_B_c_390_n N_B_c_391_n Vss PM_G4_MAJ3_N2_B
x_PM_G4_MAJ3_N2_C N_C_XI13.X0_S N_C_XI12.X0_S N_C_c_409_n N_C_c_422_p
+ N_C_c_410_n N_C_c_412_n C Vss PM_G4_MAJ3_N2_C
x_PM_G4_MAJ3_N2_Z N_Z_XI15.X0_D N_Z_XI13.X0_D N_Z_XI14.X0_D N_Z_XI12.X0_D
+ N_Z_c_427_n N_Z_c_451_n N_Z_c_432_n Z Vss PM_G4_MAJ3_N2_Z
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI11.X0_PGD 0.00200884f
cc_2 N_VDD_XI0.X0_PGD N_VSS_XI10.X0_PGD 0.0020057f
cc_3 N_VDD_c_3_p N_VSS_XI10.X0_PGD 2.76462e-19
cc_4 N_VDD_c_4_p N_VSS_c_81_n 0.00200884f
cc_5 N_VDD_c_5_p N_VSS_c_81_n 3.23379e-19
cc_6 N_VDD_c_6_p N_VSS_c_83_n 2.76462e-19
cc_7 N_VDD_c_5_p N_VSS_c_83_n 3.9313e-19
cc_8 N_VDD_c_8_p N_VSS_c_85_n 0.0020057f
cc_9 N_VDD_c_9_p N_VSS_c_85_n 2.84318e-19
cc_10 N_VDD_c_9_p N_VSS_c_87_n 3.9313e-19
cc_11 N_VDD_c_6_p N_VSS_c_88_n 4.35319e-19
cc_12 N_VDD_c_5_p N_VSS_c_88_n 0.00161703f
cc_13 N_VDD_c_13_p N_VSS_c_88_n 9.22325e-19
cc_14 N_VDD_c_14_p N_VSS_c_88_n 3.48267e-19
cc_15 N_VDD_c_3_p N_VSS_c_92_n 4.76491e-19
cc_16 N_VDD_c_9_p N_VSS_c_92_n 0.00161703f
cc_17 N_VDD_c_17_p N_VSS_c_92_n 8.59637e-19
cc_18 N_VDD_c_18_p N_VSS_c_92_n 3.48267e-19
cc_19 N_VDD_c_13_p N_VSS_c_96_n 8.49247e-19
cc_20 N_VDD_XI0.X0_PGD N_VSS_c_97_n 2.8629e-19
cc_21 N_VDD_c_17_p N_VSS_c_97_n 0.00515616f
cc_22 N_VDD_c_18_p N_VSS_c_97_n 9.58524e-19
cc_23 N_VDD_c_9_p N_VSS_c_100_n 0.00401341f
cc_24 N_VDD_c_6_p N_VSS_c_101_n 3.66936e-19
cc_25 N_VDD_c_5_p N_VSS_c_101_n 2.26455e-19
cc_26 N_VDD_c_13_p N_VSS_c_101_n 3.99794e-19
cc_27 N_VDD_c_14_p N_VSS_c_101_n 6.489e-19
cc_28 N_VDD_c_9_p N_VSS_c_105_n 2.26455e-19
cc_29 N_VDD_c_17_p N_VSS_c_105_n 3.99794e-19
cc_30 N_VDD_c_18_p N_VSS_c_105_n 6.489e-19
cc_31 N_VDD_c_6_p N_VSS_c_108_n 0.00335989f
cc_32 N_VDD_c_32_p N_VSS_c_108_n 0.00777551f
cc_33 N_VDD_c_3_p N_VSS_c_108_n 0.0031218f
cc_34 N_VDD_c_34_p N_VSS_c_108_n 0.00104624f
cc_35 N_VDD_c_35_p N_VSS_c_108_n 0.0010706f
cc_36 N_VDD_c_5_p N_VSS_c_113_n 0.00329944f
cc_37 N_VDD_c_37_p N_VSS_c_113_n 3.33664e-19
cc_38 N_VDD_c_38_p N_VSS_c_115_n 0.00106538f
cc_39 N_VDD_c_39_p N_VSS_c_116_n 3.33664e-19
cc_40 N_VDD_c_9_p N_VSS_c_116_n 0.00329944f
cc_41 N_VDD_c_41_p N_VSS_c_118_n 0.00106538f
cc_42 N_VDD_c_5_p N_VSS_c_119_n 0.00554732f
cc_43 N_VDD_c_5_p N_VSS_c_120_n 7.74609e-19
cc_44 N_VDD_c_9_p N_VSS_c_121_n 7.74609e-19
cc_45 N_VDD_XI0.X0_PGD N_A_c_161_n 3.94724e-19
cc_46 N_VDD_XI0.X0_PGD N_A_c_162_n 4.99274e-19
cc_47 N_VDD_c_5_p N_A_c_162_n 2.55296e-19
cc_48 N_VDD_c_9_p N_A_c_162_n 2.95925e-19
cc_49 N_VDD_c_17_p N_A_c_162_n 3.33497e-19
cc_50 N_VDD_c_18_p N_A_c_162_n 2.46105e-19
cc_51 N_VDD_c_13_p N_A_c_167_n 5.45771e-19
cc_52 N_VDD_c_14_p N_A_c_167_n 4.10732e-19
cc_53 N_VDD_c_32_p N_A_c_169_n 9.17955e-19
cc_54 N_VDD_c_32_p N_A_c_170_n 4.71221e-19
cc_55 N_VDD_c_55_p N_BI_c_239_n 3.43419e-19
cc_56 N_VDD_c_37_p N_BI_c_239_n 3.72199e-19
cc_57 N_VDD_c_55_p N_BI_c_241_n 3.48267e-19
cc_58 N_VDD_c_5_p N_BI_c_241_n 4.22613e-19
cc_59 N_VDD_c_37_p N_BI_c_241_n 5.2846e-19
cc_60 N_VDD_XI9.X0_PGD N_AI_XI15.X0_PGD 2.83823e-19
cc_61 N_VDD_XI0.X0_PGD N_AI_XI15.X0_PGD 3.10667e-19
cc_62 N_VDD_c_62_p N_AI_c_299_n 2.83823e-19
cc_63 N_VDD_c_63_p N_AI_c_300_n 3.10667e-19
cc_64 N_VDD_c_64_p N_AI_c_301_n 3.43419e-19
cc_65 N_VDD_c_39_p N_AI_c_301_n 3.72199e-19
cc_66 N_VDD_c_64_p N_AI_c_303_n 3.48267e-19
cc_67 N_VDD_c_39_p N_AI_c_303_n 5.226e-19
cc_68 N_VDD_c_9_p N_AI_c_303_n 4.34701e-19
cc_69 N_VDD_c_17_p N_AI_c_306_n 9.61607e-19
cc_70 N_VDD_XI9.X0_PGD N_B_c_341_n 3.99218e-19
cc_71 N_VDD_c_32_p N_B_c_342_n 3.87456e-19
cc_72 N_VDD_c_72_p B 3.02565e-19
cc_73 N_VDD_c_13_p B 4.44319e-19
cc_74 N_VDD_c_14_p B 3.49905e-19
cc_75 N_VDD_c_13_p N_B_c_346_n 3.43988e-19
cc_76 N_VDD_c_14_p N_B_c_346_n 2.68747e-19
cc_77 N_VDD_c_18_p N_B_c_346_n 4.88234e-19
cc_78 N_VSS_XI10.X0_PGD N_A_c_161_n 3.91527e-19
cc_79 N_VSS_c_123_p N_A_c_172_n 3.43419e-19
cc_80 N_VSS_c_123_p N_A_c_162_n 2.69869e-19
cc_81 N_VSS_c_125_p N_A_c_162_n 5.38503e-19
cc_82 N_VSS_c_96_n N_A_c_162_n 3.16844e-19
cc_83 N_VSS_c_97_n N_A_c_162_n 8.92829e-19
cc_84 N_VSS_c_100_n N_A_c_162_n 2.86582e-19
cc_85 N_VSS_c_119_n N_A_c_162_n 2.99293e-19
cc_86 N_VSS_c_96_n N_A_c_179_n 0.00223349f
cc_87 N_VSS_c_96_n N_A_c_167_n 0.00150218f
cc_88 N_VSS_c_92_n N_A_c_169_n 3.34005e-19
cc_89 N_VSS_c_105_n N_A_c_169_n 6.63553e-19
cc_90 N_VSS_c_108_n N_A_c_169_n 5.04162e-19
cc_91 N_VSS_c_135_p N_A_c_170_n 2.02217e-19
cc_92 N_VSS_c_92_n N_A_c_170_n 3.2351e-19
cc_93 N_VSS_c_105_n N_A_c_170_n 2.68747e-19
cc_94 N_VSS_c_123_p N_BI_c_239_n 3.43419e-19
cc_95 N_VSS_c_123_p N_BI_c_241_n 3.48267e-19
cc_96 N_VSS_c_96_n N_BI_c_241_n 0.00105024f
cc_97 N_VSS_c_108_n N_BI_c_241_n 9.87959e-19
cc_98 N_VSS_c_119_n N_BI_c_241_n 5.43103e-19
cc_99 N_VSS_c_96_n N_BI_c_249_n 4.76944e-19
cc_100 N_VSS_c_119_n N_BI_c_249_n 6.52328e-19
cc_101 N_VSS_c_125_p N_AI_c_301_n 3.43419e-19
cc_102 N_VSS_c_97_n N_AI_c_301_n 3.48267e-19
cc_103 N_VSS_c_125_p N_AI_c_303_n 3.48267e-19
cc_104 N_VSS_c_92_n N_AI_c_303_n 0.00173332f
cc_105 N_VSS_c_97_n N_AI_c_303_n 0.00144307f
cc_106 N_VSS_c_108_n N_AI_c_303_n 0.00107717f
cc_107 N_VSS_c_97_n N_AI_c_306_n 0.0019327f
cc_108 N_VSS_c_100_n N_AI_c_306_n 0.0067288f
cc_109 N_VSS_c_97_n N_AI_c_315_n 2.82216e-19
cc_110 N_VSS_c_100_n N_AI_c_316_n 0.00177928f
cc_111 N_VSS_XI11.X0_PGD N_B_c_341_n 3.95536e-19
cc_112 N_VSS_c_108_n N_B_c_342_n 7.63393e-19
cc_113 N_VSS_c_96_n N_B_c_351_n 5.01254e-19
cc_114 N_VSS_c_125_p N_C_c_409_n 3.43419e-19
cc_115 N_VSS_c_125_p N_C_c_410_n 3.48267e-19
cc_116 N_VSS_c_97_n N_C_c_410_n 6.01757e-19
cc_117 N_A_c_187_p N_BI_XI15.X0_CG 2.06538e-19
cc_118 N_A_XI14.X0_PGD N_BI_c_252_n 9.65637e-19
cc_119 N_A_c_162_n N_BI_c_241_n 3.93183e-19
cc_120 N_A_c_179_n N_BI_c_241_n 3.15833e-19
cc_121 N_A_c_179_n N_BI_c_249_n 0.00163472f
cc_122 N_A_c_187_p N_BI_c_249_n 8.66815e-19
cc_123 N_A_c_187_p N_BI_c_257_n 4.7863e-19
cc_124 N_A_c_179_n N_BI_c_258_n 3.37713e-19
cc_125 N_A_XI14.X0_PGD N_BI_c_259_n 0.00245019f
cc_126 N_A_c_187_p N_BI_c_260_n 0.00112715f
cc_127 N_A_c_162_n N_BI_c_261_n 7.8464e-19
cc_128 N_A_XI14.X0_PGD N_AI_XI15.X0_PGD 0.0173811f
cc_129 N_A_c_179_n N_AI_XI15.X0_PGD 7.90282e-19
cc_130 N_A_c_187_p N_AI_XI15.X0_PGD 0.00103582f
cc_131 N_A_c_201_p N_AI_c_299_n 0.00196947f
cc_132 N_A_c_187_p N_AI_c_299_n 9.91291e-19
cc_133 N_A_c_203_p N_AI_c_300_n 0.00200674f
cc_134 N_A_c_161_n N_AI_c_301_n 7.16634e-19
cc_135 N_A_c_162_n N_AI_c_303_n 8.04759e-19
cc_136 N_A_c_162_n N_AI_c_306_n 0.00148587f
cc_137 N_A_XI14.X0_PGD N_B_XI14.X0_CG 9.65637e-19
cc_138 N_A_c_161_n N_B_c_341_n 0.00297252f
cc_139 N_A_c_162_n N_B_c_341_n 5.2287e-19
cc_140 N_A_c_170_n N_B_c_355_n 4.73714e-19
cc_141 N_A_c_179_n N_B_c_342_n 5.60543e-19
cc_142 N_A_c_162_n B 0.00101165f
cc_143 N_A_c_179_n B 7.63651e-19
cc_144 N_A_c_187_p N_B_c_359_n 3.89825e-19
cc_145 N_A_c_215_p N_B_c_359_n 7.82672e-19
cc_146 N_A_c_216_p N_B_c_359_n 3.42845e-19
cc_147 N_A_c_161_n N_B_c_346_n 0.00100571f
cc_148 N_A_c_179_n N_B_c_346_n 2.04384e-19
cc_149 N_A_XI14.X0_PGD N_B_c_364_n 0.00312702f
cc_150 N_A_c_216_p N_B_c_364_n 2.56268e-19
cc_151 N_A_c_162_n N_B_c_351_n 0.00214888f
cc_152 N_A_c_179_n N_B_c_351_n 0.00203212f
cc_153 N_A_c_223_p N_B_c_351_n 3.75372e-19
cc_154 N_A_c_187_p N_B_c_351_n 5.5912e-19
cc_155 N_A_c_162_n N_B_c_370_n 4.2957e-19
cc_156 N_A_c_162_n N_B_c_371_n 2.29222e-19
cc_157 N_A_c_172_n N_Z_c_427_n 3.43419e-19
cc_158 N_A_c_228_p N_Z_c_427_n 3.43419e-19
cc_159 N_A_c_223_p N_Z_c_427_n 3.48267e-19
cc_160 N_A_c_230_p N_Z_c_427_n 3.48267e-19
cc_161 N_A_c_187_p N_Z_c_427_n 7.95142e-19
cc_162 N_A_XI14.X0_PGD N_Z_c_432_n 6.68421e-19
cc_163 N_A_c_172_n N_Z_c_432_n 3.48267e-19
cc_164 N_A_c_228_p N_Z_c_432_n 3.48267e-19
cc_165 N_A_c_179_n N_Z_c_432_n 0.00126628f
cc_166 N_A_c_223_p N_Z_c_432_n 7.9714e-19
cc_167 N_A_c_230_p N_Z_c_432_n 8.16241e-19
cc_168 N_A_c_187_p N_Z_c_432_n 0.00136994f
cc_169 N_BI_XI15.X0_CG N_AI_XI15.X0_PGD 9.47088e-19
cc_170 N_BI_c_258_n N_AI_XI15.X0_PGD 0.00312702f
cc_171 N_BI_c_261_n N_AI_c_303_n 3.29431e-19
cc_172 N_BI_c_249_n N_AI_c_306_n 3.35097e-19
cc_173 N_BI_c_239_n N_B_c_341_n 9.28554e-19
cc_174 N_BI_c_249_n N_B_c_342_n 0.00169958f
cc_175 N_BI_c_249_n N_B_c_374_n 7.4385e-19
cc_176 N_BI_c_257_n N_B_c_359_n 0.00182538f
cc_177 N_BI_c_259_n N_B_c_359_n 4.99367e-19
cc_178 N_BI_c_260_n N_B_c_359_n 0.00165504f
cc_179 N_BI_c_258_n N_B_c_378_n 0.00520211f
cc_180 N_BI_c_259_n N_B_c_378_n 7.2092e-19
cc_181 N_BI_c_257_n N_B_c_364_n 4.99367e-19
cc_182 N_BI_c_258_n N_B_c_364_n 6.22265e-19
cc_183 N_BI_c_259_n N_B_c_364_n 0.00494186f
cc_184 N_BI_c_249_n N_B_c_351_n 0.00529659f
cc_185 N_BI_c_249_n N_B_c_371_n 2.67017e-19
cc_186 N_BI_c_260_n N_B_c_371_n 0.0013533f
cc_187 N_BI_c_280_p N_B_c_371_n 0.00340518f
cc_188 N_BI_c_249_n N_B_c_387_n 4.99817e-19
cc_189 N_BI_c_260_n N_B_c_387_n 9.41136e-19
cc_190 N_BI_c_283_p N_B_c_387_n 7.35033e-19
cc_191 N_BI_c_280_p N_B_c_390_n 0.00181541f
cc_192 N_BI_c_249_n N_B_c_391_n 0.00145499f
cc_193 N_BI_c_260_n N_B_c_391_n 8.66399e-19
cc_194 N_BI_c_249_n N_C_c_412_n 0.00107247f
cc_195 N_BI_c_257_n N_C_c_412_n 0.00130194f
cc_196 N_BI_c_283_p N_C_c_412_n 3.02033e-19
cc_197 N_BI_c_249_n N_Z_c_432_n 0.00190811f
cc_198 N_BI_c_257_n N_Z_c_432_n 0.00192905f
cc_199 N_BI_c_258_n N_Z_c_432_n 8.66889e-19
cc_200 N_BI_c_259_n N_Z_c_432_n 8.66889e-19
cc_201 N_BI_c_260_n N_Z_c_432_n 0.00107118f
cc_202 N_BI_c_280_p N_Z_c_432_n 0.00210701f
cc_203 N_BI_c_283_p N_Z_c_432_n 0.00100479f
cc_204 N_AI_XI15.X0_PGD N_B_c_393_n 9.65637e-19
cc_205 N_AI_c_306_n N_B_c_374_n 4.95395e-19
cc_206 N_AI_c_315_n N_B_c_374_n 3.42845e-19
cc_207 N_AI_XI15.X0_PGD N_B_c_378_n 0.00312702f
cc_208 N_AI_c_315_n N_B_c_378_n 2.56268e-19
cc_209 N_AI_c_306_n N_B_c_351_n 0.00314548f
cc_210 N_AI_c_306_n N_B_c_370_n 2.5452e-19
cc_211 N_AI_c_306_n N_B_c_371_n 2.35352e-19
cc_212 N_AI_c_306_n N_C_c_410_n 0.00152957f
cc_213 N_AI_c_306_n N_C_c_412_n 0.0018056f
cc_214 N_AI_XI15.X0_PGD N_Z_c_432_n 3.73496e-19
cc_215 N_B_c_351_n N_C_c_410_n 5.20324e-19
cc_216 N_B_c_359_n N_C_c_412_n 9.16187e-19
cc_217 N_B_c_351_n N_C_c_412_n 3.71107e-19
cc_218 N_B_c_387_n N_C_c_412_n 0.00455868f
cc_219 N_B_c_374_n N_Z_c_432_n 0.00210508f
cc_220 N_B_c_359_n N_Z_c_432_n 0.0019232f
cc_221 N_B_c_364_n N_Z_c_432_n 8.66889e-19
cc_222 N_B_c_371_n N_Z_c_432_n 4.75654e-19
cc_223 N_C_c_409_n N_Z_c_451_n 3.43419e-19
cc_224 N_C_c_422_p N_Z_c_451_n 3.43419e-19
cc_225 N_C_c_410_n N_Z_c_451_n 3.48267e-19
cc_226 N_C_c_412_n N_Z_c_451_n 3.48267e-19
cc_227 N_C_c_410_n N_Z_c_432_n 6.20216e-19
cc_228 N_C_c_412_n N_Z_c_432_n 0.00126042f
*
.ends
*
*
.subckt MAJ3_HPNW8 A B C Y VDD VSS
xgate (VDD VSS A B C Y) G4_MAJ3_N2
.ends
*
* File: G3_MIN3_T6_N2.pex.netlist
* Created: Fri Apr  1 16:54:39 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MIN3_T6_N2_VSS 2 4 6 8 10 12 27 32 37 40 42 45 53 57 60 65 70 75
+ 88 89 93 99 101 106 109 Vss
c66 107 Vss 6.43136e-19
c67 106 Vss 0.0038619f
c68 101 Vss 0.00207473f
c69 99 Vss 0.0082602f
c70 94 Vss 0.00137551f
c71 93 Vss 0.00772839f
c72 89 Vss 6.57551e-19
c73 88 Vss 0.00490261f
c74 75 Vss 0.00537019f
c75 70 Vss 7.10513e-22
c76 65 Vss 0.00231683f
c77 60 Vss 0.00177007f
c78 57 Vss 0.00552514f
c79 53 Vss 0.00488234f
c80 45 Vss 0.0850774f
c81 42 Vss 0.0849587f
c82 37 Vss 0.0679309f
c83 32 Vss 0.103906f
c84 27 Vss 0.307039f
c85 22 Vss 0.141189f
c86 10 Vss 0.134855f
c87 8 Vss 0.00171956f
c88 6 Vss 0.135276f
c89 2 Vss 0.134005f
r90 106 109 0.326018
r91 105 106 4.58464
r92 101 105 0.655813
r93 100 107 0.494161
r94 99 109 0.326018
r95 99 100 13.0037
r96 95 107 0.128424
r97 93 107 0.494161
r98 93 94 10.0862
r99 88 94 0.652036
r100 87 89 0.655813
r101 87 88 12.7536
r102 70 101 1.82344
r103 65 95 5.2515
r104 60 75 1.16709
r105 60 89 1.82344
r106 57 70 1.16709
r107 53 65 1.16709
r108 45 47 1.8672
r109 42 44 1.8672
r110 40 75 0.50025
r111 37 40 1.92555
r112 33 47 0.0685365
r113 32 34 0.652036
r114 32 33 2.8008
r115 29 47 0.5835
r116 28 42 0.0685365
r117 27 45 0.0685365
r118 27 28 10.9698
r119 24 44 0.5835
r120 23 37 0.0685365
r121 22 44 0.0685365
r122 22 23 4.7847
r123 12 57 0.185659
r124 10 34 3.8511
r125 8 53 0.185659
r126 6 29 3.8511
r127 4 53 0.185659
r128 2 24 3.8511
.ends

.subckt PM_G3_MIN3_T6_N2_VDD 2 4 6 8 10 12 27 32 42 45 53 57 60 61 63 65 69 71
+ 73 78 81 83 Vss
c76 83 Vss 0.00671487f
c77 79 Vss 7.78098e-19
c78 78 Vss 0.00468194f
c79 73 Vss 0.00129457f
c80 71 Vss 0.0122041f
c81 69 Vss 0.00238015f
c82 65 Vss 0.00185683f
c83 63 Vss 7.50392e-19
c84 62 Vss 0.0017907f
c85 61 Vss 0.007913f
c86 60 Vss 0.00707888f
c87 57 Vss 0.00500133f
c88 53 Vss 0.00483876f
c89 45 Vss 0.0849087f
c90 42 Vss 0.0854801f
c91 38 Vss 0.0711342f
c92 32 Vss 0.106714f
c93 27 Vss 0.308162f
c94 22 Vss 0.144473f
c95 12 Vss 0.13249f
c96 8 Vss 0.133305f
c97 6 Vss 0.00171956f
c98 4 Vss 0.133098f
r99 78 81 0.349767
r100 77 78 4.58464
r101 73 81 0.306046
r102 73 75 1.82344
r103 72 79 0.494161
r104 71 77 0.652036
r105 71 72 13.0037
r106 67 79 0.128424
r107 67 69 5.2515
r108 65 83 1.16709
r109 63 65 1.82344
r110 61 79 0.494161
r111 61 62 10.0862
r112 60 63 0.655813
r113 59 62 0.652036
r114 59 60 12.7536
r115 57 75 1.16709
r116 53 69 1.16709
r117 45 46 1.8672
r118 42 43 1.8672
r119 38 83 0.50025
r120 38 40 1.92555
r121 33 45 0.0685365
r122 32 34 0.652036
r123 32 33 2.8008
r124 29 45 0.5835
r125 28 43 0.0685365
r126 27 46 0.0685365
r127 27 28 10.9698
r128 24 42 0.5835
r129 23 40 0.0685365
r130 22 42 0.0685365
r131 22 23 4.7847
r132 12 34 3.8511
r133 10 57 0.185659
r134 8 29 3.8511
r135 6 53 0.185659
r136 4 24 3.8511
r137 2 53 0.185659
.ends

.subckt PM_G3_MIN3_T6_N2_Z 2 4 6 8 10 12 32 36 41 45 49 53 55 59 63 67 Vss
c60 67 Vss 3.51451e-19
c61 65 Vss 2.45386e-19
c62 63 Vss 0.00102688f
c63 59 Vss 7.58182e-19
c64 55 Vss 0.00456155f
c65 53 Vss 6.51205e-19
c66 49 Vss 6.88903e-19
c67 45 Vss 0.00781677f
c68 41 Vss 0.00689463f
c69 36 Vss 0.00387467f
c70 32 Vss 0.00319091f
c71 12 Vss 0.00171956f
c72 10 Vss 0.00171956f
r73 61 67 0.494161
r74 61 63 3.04254
r75 57 67 0.494161
r76 57 59 3.04254
r77 56 65 0.128424
r78 55 67 0.128424
r79 55 56 10.3363
r80 51 65 0.494161
r81 51 53 3.04254
r82 47 65 0.494161
r83 47 49 3.04254
r84 45 63 1.16709
r85 41 59 1.16709
r86 36 53 1.16709
r87 32 49 1.16709
r88 12 45 0.185659
r89 10 41 0.185659
r90 8 45 0.185659
r91 6 41 0.185659
r92 4 36 0.185659
r93 2 32 0.185659
.ends

.subckt PM_G3_MIN3_T6_N2_C 2 4 6 8 14 20 26 29 33 38 43 Vss
c35 43 Vss 0.00523941f
c36 38 Vss 0.00156891f
c37 33 Vss 0.00543691f
c38 29 Vss 3.56438e-22
c39 20 Vss 0.377731f
c40 14 Vss 0.380603f
r41 33 43 1.16709
r42 29 38 1.16709
r43 29 33 10.0654
r44 26 29 0.0729375
r45 20 43 0.50025
r46 14 38 0.50025
r47 6 8 10.1529
r48 6 20 3.09255
r49 2 4 10.1529
r50 2 14 3.09255
.ends

.subckt PM_G3_MIN3_T6_N2_B 2 4 6 8 17 18 26 29 35 Vss
c31 35 Vss 0.00144085f
c32 26 Vss 0.0839596f
c33 18 Vss 0.0346166f
c34 17 Vss 0.0963518f
c35 6 Vss 0.399392f
c36 2 Vss 0.447969f
r37 32 35 1.16709
r38 29 32 0.0833571
r39 24 35 0.0476429
r40 24 26 1.92555
r41 17 19 0.652036
r42 17 18 2.8008
r43 14 26 0.0685365
r44 13 18 0.652036
r45 6 8 10.1529
r46 6 19 3.8511
r47 4 14 3.8511
r48 2 4 10.1529
r49 2 13 3.8511
.ends

.subckt PM_G3_MIN3_T6_N2_A 2 4 6 8 17 29 34 38 41 46 Vss
c28 46 Vss 0.00532741f
c29 41 Vss 0.00134116f
c30 34 Vss 0.00178881f
c31 26 Vss 0.0871242f
c32 6 Vss 0.406031f
c33 2 Vss 0.376065f
r34 34 46 1.16709
r35 34 38 0.0416786
r36 29 41 1.16709
r37 29 34 5.03269
r38 24 46 0.0476429
r39 24 26 1.92555
r40 19 26 0.0685365
r41 17 41 0.50025
r42 8 19 3.8511
r43 6 8 10.1529
r44 4 17 3.09255
r45 2 4 10.1529
.ends

.subckt G3_MIN3_T6_N2  VSS VDD Z C B A
*
* A	A
* B	B
* C	C
* Z	Z
* VDD	VDD
* VSS	VSS
XI17.X0 N_Z_XI17.X0_D N_VSS_XI17.X0_PGD N_C_XI17.X0_CG N_B_XI17.X0_PGS
+ N_VDD_XI17.X0_S TIGFET_HPNW8
XI14.X0 N_Z_XI14.X0_D N_VDD_XI14.X0_PGD N_C_XI14.X0_CG N_B_XI14.X0_PGS
+ N_VSS_XI14.X0_S TIGFET_HPNW8
XI19.X0 N_Z_XI19.X0_D N_VSS_XI19.X0_PGD N_A_XI19.X0_CG N_B_XI19.X0_PGS
+ N_VDD_XI19.X0_S TIGFET_HPNW8
XI16.X0 N_Z_XI16.X0_D N_VDD_XI16.X0_PGD N_A_XI16.X0_CG N_B_XI16.X0_PGS
+ N_VSS_XI16.X0_S TIGFET_HPNW8
XI18.X0 N_Z_XI18.X0_D N_VSS_XI18.X0_PGD N_C_XI18.X0_CG N_A_XI18.X0_PGS
+ N_VDD_XI18.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_VDD_XI15.X0_PGD N_C_XI15.X0_CG N_A_XI15.X0_PGS
+ N_VSS_XI15.X0_S TIGFET_HPNW8
*
x_PM_G3_MIN3_T6_N2_VSS N_VSS_XI17.X0_PGD N_VSS_XI14.X0_S N_VSS_XI19.X0_PGD
+ N_VSS_XI16.X0_S N_VSS_XI18.X0_PGD N_VSS_XI15.X0_S N_VSS_c_19_p N_VSS_c_21_p
+ N_VSS_c_7_p N_VSS_c_13_p N_VSS_c_14_p N_VSS_c_50_p N_VSS_c_4_p N_VSS_c_22_p
+ N_VSS_c_8_p N_VSS_c_28_p N_VSS_c_6_p N_VSS_c_9_p N_VSS_c_10_p N_VSS_c_11_p
+ N_VSS_c_18_p N_VSS_c_47_p N_VSS_c_24_p N_VSS_c_66_p VSS Vss
+ PM_G3_MIN3_T6_N2_VSS
x_PM_G3_MIN3_T6_N2_VDD N_VDD_XI17.X0_S N_VDD_XI14.X0_PGD N_VDD_XI19.X0_S
+ N_VDD_XI16.X0_PGD N_VDD_XI18.X0_S N_VDD_XI15.X0_PGD N_VDD_c_70_n N_VDD_c_141_p
+ N_VDD_c_134_p N_VDD_c_133_p N_VDD_c_71_n N_VDD_c_72_n N_VDD_c_73_n
+ N_VDD_c_78_n N_VDD_c_82_n N_VDD_c_83_n N_VDD_c_85_n N_VDD_c_86_n N_VDD_c_88_n
+ N_VDD_c_123_p VDD N_VDD_c_91_n Vss PM_G3_MIN3_T6_N2_VDD
x_PM_G3_MIN3_T6_N2_Z N_Z_XI17.X0_D N_Z_XI14.X0_D N_Z_XI19.X0_D N_Z_XI16.X0_D
+ N_Z_XI18.X0_D N_Z_XI15.X0_D N_Z_c_143_n N_Z_c_144_n N_Z_c_166_n N_Z_c_146_n
+ N_Z_c_150_n N_Z_c_152_n N_Z_c_155_n N_Z_c_180_n N_Z_c_157_n Z Vss
+ PM_G3_MIN3_T6_N2_Z
x_PM_G3_MIN3_T6_N2_C N_C_XI17.X0_CG N_C_XI14.X0_CG N_C_XI18.X0_CG N_C_XI15.X0_CG
+ N_C_c_203_n N_C_c_204_n C N_C_c_210_n N_C_c_205_n N_C_c_207_n N_C_c_208_n Vss
+ PM_G3_MIN3_T6_N2_C
x_PM_G3_MIN3_T6_N2_B N_B_XI17.X0_PGS N_B_XI14.X0_PGS N_B_XI19.X0_PGS
+ N_B_XI16.X0_PGS N_B_c_242_n N_B_c_243_n N_B_c_251_n B N_B_c_253_n Vss
+ PM_G3_MIN3_T6_N2_B
x_PM_G3_MIN3_T6_N2_A N_A_XI19.X0_CG N_A_XI16.X0_CG N_A_XI18.X0_PGS
+ N_A_XI15.X0_PGS N_A_c_283_n N_A_c_270_n N_A_c_272_n A N_A_c_278_n N_A_c_279_n
+ Vss PM_G3_MIN3_T6_N2_A
cc_1 N_VSS_XI17.X0_PGD N_VDD_XI14.X0_PGD 6.38995e-19
cc_2 N_VSS_XI19.X0_PGD N_VDD_XI16.X0_PGD 6.38995e-19
cc_3 N_VSS_XI18.X0_PGD N_VDD_XI15.X0_PGD 6.25013e-19
cc_4 N_VSS_c_4_p N_VDD_c_70_n 4.60829e-19
cc_5 N_VSS_c_4_p N_VDD_c_71_n 8.28334e-19
cc_6 N_VSS_c_6_p N_VDD_c_72_n 2.52506e-19
cc_7 N_VSS_c_7_p N_VDD_c_73_n 2.61781e-19
cc_8 N_VSS_c_8_p N_VDD_c_73_n 0.00161042f
cc_9 N_VSS_c_9_p N_VDD_c_73_n 0.00119047f
cc_10 N_VSS_c_10_p N_VDD_c_73_n 0.00515748f
cc_11 N_VSS_c_11_p N_VDD_c_73_n 0.00184852f
cc_12 N_VSS_c_7_p N_VDD_c_78_n 8.70611e-19
cc_13 N_VSS_c_13_p N_VDD_c_78_n 3.72495e-19
cc_14 N_VSS_c_14_p N_VDD_c_78_n 7.57734e-19
cc_15 N_VSS_c_8_p N_VDD_c_78_n 9.95408e-19
cc_16 N_VSS_c_10_p N_VDD_c_82_n 0.00175335f
cc_17 N_VSS_c_8_p N_VDD_c_83_n 5.25611e-19
cc_18 N_VSS_c_18_p N_VDD_c_83_n 4.37902e-19
cc_19 N_VSS_c_19_p N_VDD_c_85_n 0.00120274f
cc_20 N_VSS_c_19_p N_VDD_c_86_n 8.56547e-19
cc_21 N_VSS_c_21_p N_VDD_c_86_n 8.4058e-19
cc_22 N_VSS_c_22_p N_VDD_c_88_n 2.52506e-19
cc_23 N_VSS_c_6_p N_VDD_c_88_n 3.68696e-19
cc_24 N_VSS_c_24_p N_VDD_c_88_n 0.0014668f
cc_25 N_VSS_c_9_p N_VDD_c_91_n 5.6037e-19
cc_26 N_VSS_c_9_p N_Z_c_143_n 0.00379015f
cc_27 N_VSS_c_4_p N_Z_c_144_n 3.43419e-19
cc_28 N_VSS_c_28_p N_Z_c_144_n 3.48267e-19
cc_29 N_VSS_c_4_p N_Z_c_146_n 3.43419e-19
cc_30 N_VSS_c_22_p N_Z_c_146_n 3.43419e-19
cc_31 N_VSS_c_28_p N_Z_c_146_n 3.48267e-19
cc_32 N_VSS_c_6_p N_Z_c_146_n 3.48267e-19
cc_33 N_VSS_c_8_p N_Z_c_150_n 6.97647e-19
cc_34 N_VSS_c_10_p N_Z_c_150_n 0.00155764f
cc_35 N_VSS_c_4_p N_Z_c_152_n 3.48267e-19
cc_36 N_VSS_c_28_p N_Z_c_152_n 5.03066e-19
cc_37 N_VSS_c_18_p N_Z_c_152_n 5.19985e-19
cc_38 N_VSS_c_28_p N_Z_c_155_n 9.68887e-19
cc_39 N_VSS_c_18_p N_Z_c_155_n 2.48288e-19
cc_40 N_VSS_c_4_p N_Z_c_157_n 3.48267e-19
cc_41 N_VSS_c_22_p N_Z_c_157_n 3.48267e-19
cc_42 N_VSS_c_28_p N_Z_c_157_n 4.99861e-19
cc_43 N_VSS_c_6_p N_Z_c_157_n 5.71987e-19
cc_44 N_VSS_XI17.X0_PGD N_C_c_203_n 4.30517e-19
cc_45 N_VSS_XI18.X0_PGD N_C_c_204_n 5.02359e-19
cc_46 N_VSS_c_18_p N_C_c_205_n 2.62126e-19
cc_47 N_VSS_c_47_p N_C_c_205_n 5.86314e-19
cc_48 N_VSS_XI17.X0_PGD N_C_c_207_n 4.3583e-19
cc_49 N_VSS_XI18.X0_PGD N_C_c_208_n 3.76133e-19
cc_50 N_VSS_c_50_p N_C_c_208_n 2.17009e-19
cc_51 N_VSS_XI17.X0_PGD N_B_XI17.X0_PGS 0.00109504f
cc_52 N_VSS_XI19.X0_PGD N_B_XI17.X0_PGS 2.15671e-19
cc_53 N_VSS_XI19.X0_PGD N_B_XI19.X0_PGS 0.00177732f
cc_54 N_VSS_XI18.X0_PGD N_B_XI19.X0_PGS 2.22194e-19
cc_55 N_VSS_c_50_p N_B_c_242_n 0.00177732f
cc_56 N_VSS_c_19_p N_B_c_243_n 0.00719168f
cc_57 N_VSS_c_14_p N_B_c_243_n 0.00109504f
cc_58 N_VSS_c_28_p B 2.11465e-19
cc_59 N_VSS_c_10_p B 2.74582e-19
cc_60 N_VSS_c_18_p B 3.96756e-19
cc_61 N_VSS_c_19_p N_A_XI19.X0_CG 2.63627e-19
cc_62 N_VSS_c_28_p N_A_c_270_n 3.13396e-19
cc_63 N_VSS_c_47_p N_A_c_270_n 5.88825e-19
cc_64 N_VSS_c_28_p N_A_c_272_n 0.00159318f
cc_65 N_VSS_c_47_p N_A_c_272_n 0.00984051f
cc_66 N_VSS_c_66_p N_A_c_272_n 0.00110288f
cc_67 N_VDD_c_71_n N_Z_c_143_n 3.43419e-19
cc_68 N_VDD_c_73_n N_Z_c_143_n 3.70842e-19
cc_69 N_VDD_c_78_n N_Z_c_143_n 3.4118e-19
cc_70 N_VDD_c_85_n N_Z_c_143_n 3.48267e-19
cc_71 N_VDD_c_91_n N_Z_c_144_n 0.00379015f
cc_72 N_VDD_c_71_n N_Z_c_166_n 3.43419e-19
cc_73 N_VDD_c_72_n N_Z_c_166_n 3.43419e-19
cc_74 N_VDD_c_85_n N_Z_c_166_n 3.48267e-19
cc_75 N_VDD_c_86_n N_Z_c_166_n 3.4118e-19
cc_76 N_VDD_c_88_n N_Z_c_166_n 3.72199e-19
cc_77 N_VDD_c_71_n N_Z_c_150_n 3.48267e-19
cc_78 N_VDD_c_73_n N_Z_c_150_n 0.00302769f
cc_79 N_VDD_c_78_n N_Z_c_150_n 6.28868e-19
cc_80 N_VDD_c_85_n N_Z_c_150_n 7.10279e-19
cc_81 N_VDD_c_83_n N_Z_c_152_n 5.83135e-19
cc_82 N_VDD_c_71_n N_Z_c_155_n 6.44146e-19
cc_83 N_VDD_c_78_n N_Z_c_155_n 2.8517e-19
cc_84 N_VDD_c_85_n N_Z_c_155_n 0.00109243f
cc_85 N_VDD_c_86_n N_Z_c_155_n 5.3605e-19
cc_86 N_VDD_c_71_n N_Z_c_180_n 3.48267e-19
cc_87 N_VDD_c_72_n N_Z_c_180_n 3.48267e-19
cc_88 N_VDD_c_85_n N_Z_c_180_n 7.22734e-19
cc_89 N_VDD_c_86_n N_Z_c_180_n 4.75018e-19
cc_90 N_VDD_c_88_n N_Z_c_180_n 8.5731e-19
cc_91 N_VDD_c_73_n N_C_c_210_n 2.63478e-19
cc_92 N_VDD_c_78_n N_C_c_210_n 0.00145322f
cc_93 N_VDD_c_85_n N_C_c_210_n 0.00137559f
cc_94 N_VDD_c_73_n N_C_c_205_n 2.14517e-19
cc_95 N_VDD_c_78_n N_C_c_205_n 7.60337e-19
cc_96 N_VDD_c_85_n N_C_c_205_n 0.00216983f
cc_97 N_VDD_c_86_n N_C_c_205_n 0.00534093f
cc_98 N_VDD_c_123_p N_C_c_205_n 7.91462e-19
cc_99 N_VDD_c_78_n N_C_c_207_n 7.51813e-19
cc_100 N_VDD_c_85_n N_C_c_207_n 8.66889e-19
cc_101 N_VDD_c_85_n N_C_c_208_n 2.22969e-19
cc_102 N_VDD_c_86_n N_C_c_208_n 2.63125e-19
cc_103 N_VDD_c_123_p N_C_c_208_n 4.2857e-19
cc_104 N_VDD_XI14.X0_PGD N_B_XI17.X0_PGS 0.00135245f
cc_105 N_VDD_XI16.X0_PGD N_B_XI17.X0_PGS 4.12959e-19
cc_106 N_VDD_c_70_n N_B_XI19.X0_PGS 0.00107949f
cc_107 N_VDD_c_70_n N_B_c_251_n 0.00255555f
cc_108 N_VDD_c_133_p N_B_c_251_n 4.12959e-19
cc_109 N_VDD_c_134_p N_B_c_253_n 0.00495207f
cc_110 N_VDD_c_91_n N_B_c_253_n 4.60491e-19
cc_111 N_VDD_XI16.X0_PGD N_A_XI19.X0_CG 4.83278e-19
cc_112 N_VDD_XI15.X0_PGD N_A_XI18.X0_PGS 0.00150004f
cc_113 N_VDD_c_86_n N_A_XI18.X0_PGS 2.04873e-19
cc_114 N_VDD_XI16.X0_PGD N_A_c_278_n 5.50272e-19
cc_115 N_VDD_XI15.X0_PGD N_A_c_279_n 3.23173e-19
cc_116 N_VDD_c_141_p N_A_c_279_n 0.00145458f
cc_117 N_VDD_c_133_p N_A_c_279_n 2.17009e-19
cc_118 N_Z_c_150_n N_C_c_203_n 2.87038e-19
cc_119 N_Z_c_152_n N_C_c_203_n 2.87038e-19
cc_120 N_Z_c_155_n N_C_c_203_n 6.35192e-19
cc_121 N_Z_c_180_n N_C_c_204_n 0.00103972f
cc_122 N_Z_c_155_n N_C_c_210_n 3.21572e-19
cc_123 N_Z_c_155_n N_C_c_205_n 0.00152991f
cc_124 N_Z_c_180_n N_C_c_205_n 2.21606e-19
cc_125 N_Z_c_155_n N_C_c_207_n 5.52863e-19
cc_126 N_Z_c_155_n N_B_XI17.X0_PGS 7.14549e-19
cc_127 N_Z_c_155_n N_B_XI19.X0_PGS 7.57192e-19
cc_128 N_Z_c_155_n B 4.22756e-19
cc_129 N_Z_c_155_n N_B_c_253_n 5.52863e-19
cc_130 N_Z_c_155_n N_A_XI19.X0_CG 6.53623e-19
cc_131 N_Z_c_155_n N_A_c_283_n 2.7527e-19
cc_132 N_Z_c_155_n N_A_c_270_n 3.25192e-19
cc_133 N_Z_c_155_n N_A_c_272_n 2.57254e-19
cc_134 N_Z_c_157_n N_A_c_272_n 4.03022e-19
cc_135 N_Z_c_155_n N_A_c_278_n 2.77593e-19
cc_136 N_C_c_203_n N_B_XI17.X0_PGS 0.00849032f
cc_137 N_C_c_207_n N_B_XI17.X0_PGS 3.76133e-19
cc_138 N_C_c_203_n N_B_XI19.X0_PGS 6.67601e-19
cc_139 N_C_c_204_n N_B_XI19.X0_PGS 4.29907e-19
cc_140 N_C_c_204_n N_A_XI19.X0_CG 0.00200107f
cc_141 N_C_c_204_n N_A_XI18.X0_PGS 0.00801113f
cc_142 N_C_c_205_n N_A_c_272_n 0.00154898f
cc_143 N_B_XI17.X0_PGS N_A_XI19.X0_CG 8.40291e-19
cc_144 N_B_XI19.X0_PGS N_A_XI19.X0_CG 0.00774979f
cc_145 B N_A_c_270_n 3.39698e-19
cc_146 N_B_c_253_n N_A_c_270_n 3.48267e-19
cc_147 B N_A_c_278_n 3.48267e-19
cc_148 N_B_c_253_n N_A_c_278_n 5.15124e-19
*
.ends
*
*
.subckt MIN3_HPNW8 A B C Y VDD VSS
xgate (VSS VDD Y C B A) G3_MIN3_T6_N2
.ends
*
* File: G4_MUX2_N2.pex.netlist
* Created: Tue Mar 15 11:14:18 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MUX2_N2_VDD 2 4 6 8 10 12 14 16 18 20 38 49 51 58 64 72 77 81 84
+ 85 89 93 95 96 99 101 105 107 111 113 115 120 122 124 125 126 127 128 134 139
+ 148 Vss
c133 148 Vss 0.00699273f
c134 139 Vss 0.00445774f
c135 134 Vss 0.00494975f
c136 128 Vss 4.52364e-19
c137 127 Vss 2.39889e-19
c138 126 Vss 4.2334e-19
c139 125 Vss 2.39889e-19
c140 122 Vss 0.00207203f
c141 120 Vss 0.00831709f
c142 115 Vss 0.00192f
c143 113 Vss 0.00621353f
c144 111 Vss 7.23227e-19
c145 107 Vss 0.00783849f
c146 105 Vss 0.0013925f
c147 101 Vss 0.00172494f
c148 99 Vss 3.98903e-19
c149 96 Vss 6.1175e-19
c150 95 Vss 0.00348383f
c151 93 Vss 0.00103115f
c152 89 Vss 0.0016395f
c153 86 Vss 0.00175544f
c154 85 Vss 0.00656595f
c155 84 Vss 0.0047574f
c156 81 Vss 0.00425172f
c157 77 Vss 0.00710807f
c158 72 Vss 0.00394783f
c159 64 Vss 9.76046e-20
c160 59 Vss 0.0805856f
c161 58 Vss 0.104002f
c162 51 Vss 1.36639e-19
c163 49 Vss 0.035607f
c164 48 Vss 0.101298f
c165 39 Vss 0.0367217f
c166 38 Vss 0.101451f
c167 18 Vss 0.134291f
c168 16 Vss 0.00143442f
c169 14 Vss 0.136641f
c170 10 Vss 0.134979f
c171 8 Vss 0.134694f
c172 6 Vss 0.136393f
c173 4 Vss 0.134706f
r174 121 128 0.551426
r175 121 122 4.58464
r176 120 128 0.551426
r177 119 120 15.5878
r178 115 128 0.0828784
r179 115 117 1.82344
r180 114 127 0.494161
r181 113 119 0.652036
r182 113 114 10.1279
r183 111 148 1.16709
r184 109 127 0.128424
r185 109 111 2.16729
r186 108 126 0.494161
r187 107 122 0.652036
r188 107 108 13.0037
r189 103 126 0.128424
r190 103 105 5.2515
r191 102 125 0.494161
r192 101 127 0.494161
r193 101 102 4.58464
r194 99 139 1.16709
r195 97 125 0.128424
r196 97 99 2.16729
r197 95 126 0.494161
r198 95 96 7.46046
r199 93 134 1.16709
r200 91 96 0.652036
r201 91 93 2.16729
r202 87 124 0.306046
r203 87 89 1.82344
r204 85 125 0.494161
r205 85 86 10.1279
r206 84 124 0.349767
r207 83 86 0.652036
r208 83 84 4.58464
r209 81 117 1.16709
r210 77 105 1.16709
r211 72 89 1.16709
r212 64 148 0.0476429
r213 64 66 1.92555
r214 59 66 0.5835
r215 58 60 0.652036
r216 58 59 2.8008
r217 55 66 0.0685365
r218 51 139 0.0476429
r219 49 51 1.45875
r220 48 52 0.652036
r221 48 51 1.45875
r222 45 49 0.652036
r223 41 134 0.0476429
r224 39 41 1.45875
r225 38 42 0.652036
r226 38 41 1.45875
r227 35 39 0.652036
r228 20 81 0.185659
r229 18 60 3.8511
r230 16 77 0.185659
r231 14 55 3.8511
r232 12 77 0.185659
r233 10 52 3.8511
r234 8 45 3.8511
r235 6 35 3.8511
r236 4 42 3.8511
r237 2 72 0.185659
.ends

.subckt PM_G4_MUX2_N2_VSS 2 4 6 8 10 12 14 16 18 20 38 39 41 48 49 59 72 77 81
+ 84 89 94 99 104 109 118 123 132 141 142 146 152 153 158 164 170 172 177 179
+ 181 182 183 184 185 Vss
c128 185 Vss 4.28045e-19
c129 184 Vss 3.62111e-19
c130 183 Vss 3.88979e-19
c131 182 Vss 3.21876e-19
c132 179 Vss 0.00491274f
c133 177 Vss 0.00148831f
c134 172 Vss 0.00130997f
c135 170 Vss 0.0025874f
c136 164 Vss 0.00591751f
c137 158 Vss 0.00396568f
c138 153 Vss 5.94991e-19
c139 152 Vss 0.00255814f
c140 146 Vss 0.00513861f
c141 142 Vss 0.00102564f
c142 141 Vss 0.00403723f
c143 132 Vss 0.00811196f
c144 123 Vss 0.00369111f
c145 118 Vss 0.00399678f
c146 109 Vss 4.35064e-19
c147 104 Vss 0.00132832f
c148 99 Vss 0.00135757f
c149 94 Vss 4.3806e-19
c150 89 Vss 9.57033e-19
c151 84 Vss 0.00151444f
c152 81 Vss 0.00400382f
c153 77 Vss 0.00617013f
c154 72 Vss 0.00549529f
c155 65 Vss 0.0783825f
c156 59 Vss 0.0350566f
c157 58 Vss 0.0688416f
c158 49 Vss 0.0347733f
c159 48 Vss 0.100344f
c160 41 Vss 9.8832e-20
c161 39 Vss 0.0350852f
c162 38 Vss 0.0994129f
c163 20 Vss 0.135394f
c164 16 Vss 0.134482f
c165 14 Vss 0.00143442f
c166 12 Vss 0.134697f
c167 10 Vss 0.135146f
c168 4 Vss 0.134814f
c169 2 Vss 0.13402f
r170 178 185 0.551426
r171 178 179 15.5878
r172 177 185 0.551426
r173 176 177 4.58464
r174 172 185 0.0828784
r175 171 184 0.494161
r176 170 179 0.652036
r177 170 171 4.41793
r178 166 184 0.128424
r179 165 183 0.494161
r180 164 176 0.652036
r181 164 165 13.0037
r182 160 183 0.128424
r183 159 182 0.494161
r184 158 184 0.494161
r185 158 159 10.2946
r186 154 182 0.128424
r187 152 183 0.494161
r188 152 153 7.46046
r189 148 153 0.652036
r190 147 181 0.326018
r191 146 182 0.494161
r192 146 147 10.1279
r193 141 181 0.326018
r194 140 142 0.655813
r195 140 141 4.58464
r196 109 172 1.82344
r197 104 132 1.16709
r198 104 166 2.16729
r199 99 160 5.2515
r200 94 123 1.16709
r201 94 154 2.16729
r202 89 118 1.16709
r203 89 148 2.16729
r204 84 142 1.82344
r205 81 109 1.16709
r206 77 99 1.16709
r207 72 84 1.16709
r208 65 132 0.0476429
r209 63 65 1.8672
r210 60 63 0.0685365
r211 58 63 0.5835
r212 58 59 2.8008
r213 55 59 0.652036
r214 51 123 0.0476429
r215 49 51 1.45875
r216 48 52 0.652036
r217 48 51 1.45875
r218 45 49 0.652036
r219 41 118 0.0476429
r220 39 41 1.45875
r221 38 42 0.652036
r222 38 41 1.45875
r223 35 39 0.652036
r224 20 60 3.8511
r225 18 81 0.185659
r226 16 55 3.8511
r227 14 77 0.185659
r228 12 52 3.8511
r229 10 45 3.8511
r230 8 77 0.185659
r231 6 72 0.185659
r232 4 35 3.8511
r233 2 42 3.8511
.ends

.subckt PM_G4_MUX2_N2_ZI 2 4 6 8 10 12 27 28 43 47 50 55 60 65 81 82 91 Vss
c67 82 Vss 9.49146e-19
c68 81 Vss 0.00328207f
c69 65 Vss 0.00492924f
c70 60 Vss 0.00114673f
c71 55 Vss 0.00119934f
c72 50 Vss 0.00186152f
c73 47 Vss 0.00662602f
c74 43 Vss 0.00662602f
c75 28 Vss 0.204565f
c76 27 Vss 9.8832e-20
c77 23 Vss 0.0247918f
c78 12 Vss 0.00143442f
c79 10 Vss 0.00143442f
c80 4 Vss 0.134965f
c81 2 Vss 0.126125f
r82 87 91 0.494161
r83 83 91 0.494161
r84 81 91 0.128424
r85 81 82 13.2121
r86 77 82 0.652036
r87 60 87 4.58464
r88 55 83 5.2515
r89 50 65 1.16709
r90 50 77 2.16729
r91 47 60 1.16709
r92 43 55 1.16709
r93 31 65 0.0476429
r94 29 31 0.326018
r95 29 31 0.1167
r96 28 32 0.652036
r97 28 31 6.7686
r98 27 65 0.357321
r99 23 31 0.326018
r100 23 27 0.40845
r101 12 47 0.185659
r102 10 43 0.185659
r103 8 47 0.185659
r104 6 43 0.185659
r105 4 32 3.8511
r106 2 27 3.44265
.ends

.subckt PM_G4_MUX2_N2_Z 2 4 13 16 19 Vss
c13 16 Vss 2.38782e-19
c14 13 Vss 0.00448964f
c15 4 Vss 0.00143442f
r16 16 19 0.0416786
r17 13 16 1.16709
r18 4 13 0.185659
r19 2 13 0.185659
.ends

.subckt PM_G4_MUX2_N2_SELI 2 4 6 8 18 21 29 33 36 38 43 44 52 57 71 76 77 Vss
c77 77 Vss 8.68628e-19
c78 76 Vss 1.71087e-19
c79 71 Vss 0.00181943f
c80 57 Vss 0.00285848f
c81 52 Vss 0.00302696f
c82 44 Vss 0.00257468f
c83 43 Vss 7.72677e-19
c84 38 Vss 0.00166363f
c85 36 Vss 3.84679e-19
c86 33 Vss 0.00302237f
c87 29 Vss 0.00550884f
c88 21 Vss 0.112078f
c89 18 Vss 1.01432e-19
c90 6 Vss 0.112115f
c91 4 Vss 0.00143442f
r92 76 77 0.655813
r93 75 76 3.501
r94 71 75 0.655813
r95 43 52 1.16709
r96 43 71 2.00578
r97 43 44 0.513084
r98 38 57 1.16709
r99 38 77 2.00578
r100 36 44 7.46046
r101 31 36 0.652036
r102 31 33 7.002
r103 29 33 1.16709
r104 21 57 0.50025
r105 18 52 0.50025
r106 8 21 3.09255
r107 6 18 3.09255
r108 4 29 0.185659
r109 2 29 0.185659
.ends

.subckt PM_G4_MUX2_N2_SEL 2 4 6 8 16 17 22 26 33 36 40 41 44 45 47 49 56 57 59
+ 64 69 Vss
c70 69 Vss 0.00270368f
c71 64 Vss 0.00315728f
c72 59 Vss 0.00270998f
c73 57 Vss 3.45787e-19
c74 56 Vss 0.00198364f
c75 49 Vss 3.06667e-19
c76 47 Vss 0.00132431f
c77 45 Vss 4.54881e-19
c78 44 Vss 0.00192809f
c79 41 Vss 0.00173298f
c80 36 Vss 9.81095e-20
c81 33 Vss 1.05421e-19
c82 26 Vss 0.112078f
c83 22 Vss 0.125771f
c84 20 Vss 0.0247918f
c85 17 Vss 0.0358516f
c86 16 Vss 0.176172f
c87 8 Vss 0.112078f
c88 2 Vss 0.139232f
r89 55 64 1.16709
r90 55 57 0.4602
r91 55 56 0.52504
r92 52 59 1.16709
r93 49 52 0.5835
r94 47 69 1.16709
r95 45 47 2.00578
r96 43 45 0.655813
r97 43 44 3.501
r98 41 44 0.655813
r99 41 57 1.49522
r100 40 56 3.04254
r101 38 49 0.0685365
r102 38 40 1.54211
r103 36 59 0.0476429
r104 33 69 0.50025
r105 26 64 0.50025
r106 22 59 0.357321
r107 20 36 0.326018
r108 20 22 0.40845
r109 17 36 6.7686
r110 16 36 0.326018
r111 16 36 0.1167
r112 13 17 0.652036
r113 8 33 3.09255
r114 6 26 3.09255
r115 4 22 3.44265
r116 2 13 3.8511
.ends

.subckt PM_G4_MUX2_N2_B 2 4 14 20 23 Vss
c30 23 Vss 0.00425113f
c31 20 Vss 3.02878e-19
c32 14 Vss 0.0853035f
c33 2 Vss 0.547212f
r34 17 23 1.16709
r35 17 20 0.0729375
r36 14 23 0.0476429
r37 11 14 1.92555
r38 7 11 0.0685365
r39 4 7 3.8511
r40 2 4 15.4044
.ends

.subckt PM_G4_MUX2_N2_A 2 4 12 14 17 23 Vss
c24 23 Vss 0.00254505f
c25 17 Vss 3.13475e-19
c26 14 Vss 0.0661045f
c27 12 Vss 1.05421e-19
c28 2 Vss 0.578847f
r29 20 23 1.16709
r30 17 20 0.0833571
r31 12 23 0.3335
r32 12 14 1.57545
r33 7 14 0.0685365
r34 2 4 15.4044
r35 2 7 4.60965
.ends

.subckt G4_MUX2_N2  VDD VSS Z SEL B A
*
* A	A
* B	B
* SEL	SEL
* Z	Z
* VSS	VSS
* VDD	VDD
XI5.X0 N_Z_XI5.X0_D N_VSS_XI5.X0_PGD N_ZI_XI5.X0_CG N_VSS_XI5.X0_PGS
+ N_VDD_XI5.X0_S TIGFET_HPNW8
XI6.X0 N_SELI_XI6.X0_D N_VDD_XI6.X0_PGD N_SEL_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VDD_XI4.X0_PGD N_ZI_XI4.X0_CG N_VDD_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW8
XI7.X0 N_SELI_XI7.X0_D N_VSS_XI7.X0_PGD N_SEL_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW8
XI11.X0 N_ZI_XI11.X0_D N_VDD_XI11.X0_PGD N_SELI_XI11.X0_CG N_B_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW8
XI9.X0 N_ZI_XI9.X0_D N_VSS_XI9.X0_PGD N_SEL_XI9.X0_CG N_B_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW8
XI10.X0 N_ZI_XI10.X0_D N_VDD_XI10.X0_PGD N_SEL_XI10.X0_CG N_A_XI10.X0_PGS
+ N_VSS_XI10.X0_S TIGFET_HPNW8
XI8.X0 N_ZI_XI8.X0_D N_VSS_XI8.X0_PGD N_SELI_XI8.X0_CG N_A_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW8
*
x_PM_G4_MUX2_N2_VDD N_VDD_XI5.X0_S N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS
+ N_VDD_XI4.X0_PGD N_VDD_XI4.X0_PGS N_VDD_XI7.X0_S N_VDD_XI11.X0_PGD
+ N_VDD_XI9.X0_S N_VDD_XI10.X0_PGD N_VDD_XI8.X0_S N_VDD_c_12_p N_VDD_c_8_p
+ N_VDD_c_115_p N_VDD_c_121_p N_VDD_c_91_p N_VDD_c_85_p N_VDD_c_15_p
+ N_VDD_c_72_p N_VDD_c_10_p N_VDD_c_9_p N_VDD_c_17_p N_VDD_c_22_p N_VDD_c_13_p
+ N_VDD_c_47_p N_VDD_c_20_p N_VDD_c_27_p N_VDD_c_5_p N_VDD_c_14_p N_VDD_c_28_p
+ N_VDD_c_16_p N_VDD_c_59_p N_VDD_c_29_p N_VDD_c_32_p VDD N_VDD_c_50_p
+ N_VDD_c_54_p N_VDD_c_57_p N_VDD_c_64_p N_VDD_c_25_p N_VDD_c_21_p N_VDD_c_100_p
+ Vss PM_G4_MUX2_N2_VDD
x_PM_G4_MUX2_N2_VSS N_VSS_XI5.X0_PGD N_VSS_XI5.X0_PGS N_VSS_XI6.X0_S
+ N_VSS_XI4.X0_S N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS N_VSS_XI11.X0_S
+ N_VSS_XI9.X0_PGD N_VSS_XI10.X0_S N_VSS_XI8.X0_PGD N_VSS_c_141_n N_VSS_c_143_n
+ N_VSS_c_202_p N_VSS_c_252_p N_VSS_c_145_n N_VSS_c_147_n N_VSS_c_227_p
+ N_VSS_c_148_n N_VSS_c_149_n N_VSS_c_150_n N_VSS_c_151_n N_VSS_c_155_n
+ N_VSS_c_159_n N_VSS_c_163_n N_VSS_c_166_n N_VSS_c_168_n N_VSS_c_171_n
+ N_VSS_c_175_n N_VSS_c_177_n N_VSS_c_178_n N_VSS_c_179_n N_VSS_c_181_n
+ N_VSS_c_184_n N_VSS_c_185_n N_VSS_c_188_n N_VSS_c_191_n N_VSS_c_192_n
+ N_VSS_c_193_n N_VSS_c_194_n VSS N_VSS_c_198_n N_VSS_c_199_n N_VSS_c_200_n
+ N_VSS_c_201_n Vss PM_G4_MUX2_N2_VSS
x_PM_G4_MUX2_N2_ZI N_ZI_XI5.X0_CG N_ZI_XI4.X0_CG N_ZI_XI11.X0_D N_ZI_XI9.X0_D
+ N_ZI_XI10.X0_D N_ZI_XI8.X0_D N_ZI_c_278_n N_ZI_c_262_n N_ZI_c_263_n
+ N_ZI_c_264_n N_ZI_c_283_n N_ZI_c_269_n N_ZI_c_271_n N_ZI_c_276_n N_ZI_c_277_n
+ N_ZI_c_298_n N_ZI_c_314_p Vss PM_G4_MUX2_N2_ZI
x_PM_G4_MUX2_N2_Z N_Z_XI5.X0_D N_Z_XI4.X0_D N_Z_c_329_n N_Z_c_332_n Z Vss
+ PM_G4_MUX2_N2_Z
x_PM_G4_MUX2_N2_SELI N_SELI_XI6.X0_D N_SELI_XI7.X0_D N_SELI_XI11.X0_CG
+ N_SELI_XI8.X0_CG N_SELI_c_342_n N_SELI_c_417_p N_SELI_c_343_n N_SELI_c_346_n
+ N_SELI_c_374_n N_SELI_c_349_n N_SELI_c_350_n N_SELI_c_352_n N_SELI_c_356_n
+ N_SELI_c_368_n N_SELI_c_370_n N_SELI_c_384_n N_SELI_c_387_n Vss
+ PM_G4_MUX2_N2_SELI
x_PM_G4_MUX2_N2_SEL N_SEL_XI6.X0_CG N_SEL_XI7.X0_CG N_SEL_XI9.X0_CG
+ N_SEL_XI10.X0_CG N_SEL_c_419_n N_SEL_c_439_n N_SEL_c_473_p N_SEL_c_474_p
+ N_SEL_c_484_p N_SEL_c_430_n SEL N_SEL_c_420_n N_SEL_c_421_n N_SEL_c_446_n
+ N_SEL_c_422_n N_SEL_c_433_n N_SEL_c_425_n N_SEL_c_462_n N_SEL_c_427_n
+ N_SEL_c_465_n N_SEL_c_428_n Vss PM_G4_MUX2_N2_SEL
x_PM_G4_MUX2_N2_B N_B_XI11.X0_PGS N_B_XI9.X0_PGS N_B_c_495_n B N_B_c_491_n Vss
+ PM_G4_MUX2_N2_B
x_PM_G4_MUX2_N2_A N_A_XI10.X0_PGS N_A_XI8.X0_PGS N_A_c_537_n N_A_c_521_n A
+ N_A_c_527_n Vss PM_G4_MUX2_N2_A
cc_1 N_VDD_XI4.X0_PGD N_VSS_XI5.X0_PGD 0.00201121f
cc_2 N_VDD_XI6.X0_PGS N_VSS_XI5.X0_PGS 2.37403e-19
cc_3 N_VDD_XI6.X0_PGD N_VSS_XI7.X0_PGD 0.00195824f
cc_4 N_VDD_XI4.X0_PGS N_VSS_XI7.X0_PGS 2.20829e-19
cc_5 N_VDD_c_5_p N_VSS_XI7.X0_PGS 2.10824e-19
cc_6 N_VDD_XI11.X0_PGD N_VSS_XI9.X0_PGD 2.24862e-19
cc_7 N_VDD_XI10.X0_PGD N_VSS_XI8.X0_PGD 2.24862e-19
cc_8 N_VDD_c_8_p N_VSS_c_141_n 0.00201121f
cc_9 N_VDD_c_9_p N_VSS_c_141_n 3.9313e-19
cc_10 N_VDD_c_10_p N_VSS_c_143_n 3.05236e-19
cc_11 N_VDD_c_9_p N_VSS_c_143_n 4.1253e-19
cc_12 N_VDD_c_12_p N_VSS_c_145_n 0.00195824f
cc_13 N_VDD_c_13_p N_VSS_c_145_n 3.03215e-19
cc_14 N_VDD_c_14_p N_VSS_c_147_n 8.80211e-19
cc_15 N_VDD_c_15_p N_VSS_c_148_n 3.1188e-19
cc_16 N_VDD_c_16_p N_VSS_c_149_n 3.4118e-19
cc_17 N_VDD_c_17_p N_VSS_c_150_n 5.69928e-19
cc_18 N_VDD_c_10_p N_VSS_c_151_n 8.67538e-19
cc_19 N_VDD_c_9_p N_VSS_c_151_n 0.00161703f
cc_20 N_VDD_c_20_p N_VSS_c_151_n 8.83788e-19
cc_21 N_VDD_c_21_p N_VSS_c_151_n 3.48267e-19
cc_22 N_VDD_c_22_p N_VSS_c_155_n 8.50587e-19
cc_23 N_VDD_c_13_p N_VSS_c_155_n 0.00161703f
cc_24 N_VDD_c_5_p N_VSS_c_155_n 0.00180638f
cc_25 N_VDD_c_25_p N_VSS_c_155_n 3.48267e-19
cc_26 N_VDD_c_20_p N_VSS_c_159_n 3.92901e-19
cc_27 N_VDD_c_27_p N_VSS_c_159_n 4.34701e-19
cc_28 N_VDD_c_28_p N_VSS_c_159_n 7.06793e-19
cc_29 N_VDD_c_29_p N_VSS_c_159_n 3.47458e-19
cc_30 N_VDD_c_5_p N_VSS_c_163_n 2.93442e-19
cc_31 N_VDD_c_14_p N_VSS_c_163_n 0.00161703f
cc_32 N_VDD_c_32_p N_VSS_c_163_n 4.28751e-19
cc_33 N_VDD_c_16_p N_VSS_c_166_n 4.19648e-19
cc_34 N_VDD_c_29_p N_VSS_c_166_n 0.00187494f
cc_35 N_VDD_c_10_p N_VSS_c_168_n 3.66936e-19
cc_36 N_VDD_c_9_p N_VSS_c_168_n 2.26455e-19
cc_37 N_VDD_c_21_p N_VSS_c_168_n 6.489e-19
cc_38 N_VDD_c_22_p N_VSS_c_171_n 3.82294e-19
cc_39 N_VDD_c_13_p N_VSS_c_171_n 2.26455e-19
cc_40 N_VDD_c_5_p N_VSS_c_171_n 9.55349e-19
cc_41 N_VDD_c_25_p N_VSS_c_171_n 6.46219e-19
cc_42 N_VDD_c_14_p N_VSS_c_175_n 2.26455e-19
cc_43 N_VDD_c_32_p N_VSS_c_175_n 3.63088e-19
cc_44 N_VDD_c_22_p N_VSS_c_177_n 3.85245e-19
cc_45 N_VDD_c_10_p N_VSS_c_178_n 4.00013e-19
cc_46 N_VDD_c_13_p N_VSS_c_179_n 0.00408997f
cc_47 N_VDD_c_47_p N_VSS_c_179_n 0.00164958f
cc_48 N_VDD_c_9_p N_VSS_c_181_n 0.0040756f
cc_49 N_VDD_c_27_p N_VSS_c_181_n 0.00132969f
cc_50 N_VDD_c_50_p N_VSS_c_181_n 0.00102696f
cc_51 N_VDD_c_9_p N_VSS_c_184_n 0.00176255f
cc_52 N_VDD_c_13_p N_VSS_c_185_n 0.00134925f
cc_53 N_VDD_c_14_p N_VSS_c_185_n 0.0059995f
cc_54 N_VDD_c_54_p N_VSS_c_185_n 0.00115121f
cc_55 N_VDD_c_27_p N_VSS_c_188_n 0.00132969f
cc_56 N_VDD_c_16_p N_VSS_c_188_n 0.00814611f
cc_57 N_VDD_c_57_p N_VSS_c_188_n 9.97418e-19
cc_58 N_VDD_c_14_p N_VSS_c_191_n 0.00456934f
cc_59 N_VDD_c_59_p N_VSS_c_192_n 4.54377e-19
cc_60 N_VDD_c_29_p N_VSS_c_193_n 0.00335336f
cc_61 N_VDD_c_5_p N_VSS_c_194_n 3.22916e-19
cc_62 N_VDD_c_29_p N_VSS_c_194_n 0.00738754f
cc_63 N_VDD_c_32_p N_VSS_c_194_n 0.00291237f
cc_64 N_VDD_c_64_p N_VSS_c_194_n 0.0010706f
cc_65 N_VDD_c_13_p N_VSS_c_198_n 7.23159e-19
cc_66 N_VDD_c_27_p N_VSS_c_199_n 0.00107375f
cc_67 N_VDD_c_14_p N_VSS_c_200_n 7.61747e-19
cc_68 N_VDD_c_29_p N_VSS_c_201_n 9.16632e-19
cc_69 N_VDD_XI4.X0_PGD N_ZI_c_262_n 3.93784e-19
cc_70 N_VDD_c_16_p N_ZI_c_263_n 3.4118e-19
cc_71 N_VDD_c_15_p N_ZI_c_264_n 3.43419e-19
cc_72 N_VDD_c_72_p N_ZI_c_264_n 3.43419e-19
cc_73 N_VDD_c_5_p N_ZI_c_264_n 3.48267e-19
cc_74 N_VDD_c_14_p N_ZI_c_264_n 3.4118e-19
cc_75 N_VDD_c_59_p N_ZI_c_264_n 3.72199e-19
cc_76 N_VDD_c_16_p N_ZI_c_269_n 3.98099e-19
cc_77 N_VDD_c_29_p N_ZI_c_269_n 7.67329e-19
cc_78 N_VDD_c_15_p N_ZI_c_271_n 3.48267e-19
cc_79 N_VDD_c_72_p N_ZI_c_271_n 3.48267e-19
cc_80 N_VDD_c_5_p N_ZI_c_271_n 4.99861e-19
cc_81 N_VDD_c_14_p N_ZI_c_271_n 3.98099e-19
cc_82 N_VDD_c_59_p N_ZI_c_271_n 5.226e-19
cc_83 N_VDD_c_25_p N_ZI_c_276_n 3.30805e-19
cc_84 N_VDD_c_13_p N_ZI_c_277_n 3.38227e-19
cc_85 N_VDD_c_85_p N_Z_c_329_n 3.43419e-19
cc_86 N_VDD_c_9_p N_Z_c_329_n 3.4118e-19
cc_87 N_VDD_c_17_p N_Z_c_329_n 3.72199e-19
cc_88 N_VDD_c_85_p N_Z_c_332_n 3.48267e-19
cc_89 N_VDD_c_9_p N_Z_c_332_n 4.58391e-19
cc_90 N_VDD_c_17_p N_Z_c_332_n 7.4527e-19
cc_91 N_VDD_c_91_p N_SELI_c_342_n 8.8401e-19
cc_92 N_VDD_c_15_p N_SELI_c_343_n 3.43419e-19
cc_93 N_VDD_c_13_p N_SELI_c_343_n 3.4118e-19
cc_94 N_VDD_c_5_p N_SELI_c_343_n 3.48267e-19
cc_95 N_VDD_c_15_p N_SELI_c_346_n 3.48267e-19
cc_96 N_VDD_c_13_p N_SELI_c_346_n 4.79144e-19
cc_97 N_VDD_c_5_p N_SELI_c_346_n 6.94315e-19
cc_98 N_VDD_c_29_p N_SELI_c_349_n 4.73641e-19
cc_99 N_VDD_c_28_p N_SELI_c_350_n 3.11429e-19
cc_100 N_VDD_c_100_p N_SELI_c_350_n 3.26631e-19
cc_101 N_VDD_XI4.X0_PGD N_SELI_c_352_n 2.33421e-19
cc_102 N_VDD_c_20_p N_SELI_c_352_n 4.24036e-19
cc_103 N_VDD_c_27_p N_SELI_c_352_n 2.6015e-19
cc_104 N_VDD_c_21_p N_SELI_c_352_n 2.91146e-19
cc_105 N_VDD_c_28_p N_SELI_c_356_n 3.43988e-19
cc_106 N_VDD_c_100_p N_SELI_c_356_n 2.68747e-19
cc_107 N_VDD_XI6.X0_PGD N_SEL_c_419_n 4.07423e-19
cc_108 N_VDD_c_14_p N_SEL_c_420_n 4.4769e-19
cc_109 N_VDD_c_29_p N_SEL_c_421_n 5.4414e-19
cc_110 N_VDD_c_14_p N_SEL_c_422_n 2.04009e-19
cc_111 N_VDD_c_16_p N_SEL_c_422_n 4.56389e-19
cc_112 N_VDD_c_29_p N_SEL_c_422_n 5.05119e-19
cc_113 N_VDD_c_15_p N_SEL_c_425_n 6.34806e-19
cc_114 N_VDD_c_5_p N_SEL_c_425_n 0.0010174f
cc_115 N_VDD_c_115_p N_SEL_c_427_n 4.97707e-19
cc_116 N_VDD_c_29_p N_SEL_c_428_n 3.66936e-19
cc_117 N_VDD_c_5_p B 0.00142218f
cc_118 N_VDD_c_14_p B 0.00141439f
cc_119 N_VDD_c_5_p N_B_c_491_n 9.67317e-19
cc_120 N_VDD_c_14_p N_B_c_491_n 0.00120343f
cc_121 N_VDD_c_121_p N_A_XI10.X0_PGS 0.00270087f
cc_122 N_VDD_c_29_p N_A_XI10.X0_PGS 0.00113883f
cc_123 N_VDD_c_16_p N_A_c_521_n 3.83429e-19
cc_124 N_VDD_c_29_p N_A_c_521_n 4.45055e-19
cc_125 N_VDD_c_28_p A 5.39847e-19
cc_126 N_VDD_c_16_p A 0.00141439f
cc_127 N_VDD_c_29_p A 4.93619e-19
cc_128 N_VDD_c_100_p A 3.48267e-19
cc_129 N_VDD_XI10.X0_PGD N_A_c_527_n 3.23173e-19
cc_130 N_VDD_c_28_p N_A_c_527_n 4.07426e-19
cc_131 N_VDD_c_16_p N_A_c_527_n 0.00124433f
cc_132 N_VDD_c_29_p N_A_c_527_n 3.66936e-19
cc_133 N_VDD_c_100_p N_A_c_527_n 6.47766e-19
cc_134 N_VSS_c_202_p N_ZI_c_278_n 9.69352e-19
cc_135 N_VSS_XI5.X0_PGD N_ZI_c_262_n 4.04227e-19
cc_136 N_VSS_c_148_n N_ZI_c_263_n 3.43419e-19
cc_137 N_VSS_c_149_n N_ZI_c_263_n 3.43419e-19
cc_138 N_VSS_c_166_n N_ZI_c_263_n 3.48267e-19
cc_139 N_VSS_c_151_n N_ZI_c_283_n 8.31001e-19
cc_140 N_VSS_c_168_n N_ZI_c_283_n 3.27324e-19
cc_141 N_VSS_c_148_n N_ZI_c_269_n 3.48267e-19
cc_142 N_VSS_c_149_n N_ZI_c_269_n 3.48267e-19
cc_143 N_VSS_c_159_n N_ZI_c_269_n 0.00100597f
cc_144 N_VSS_c_166_n N_ZI_c_269_n 4.40384e-19
cc_145 N_VSS_c_188_n N_ZI_c_269_n 4.67196e-19
cc_146 N_VSS_c_192_n N_ZI_c_269_n 6.1924e-19
cc_147 N_VSS_c_194_n N_ZI_c_269_n 0.0017026f
cc_148 N_VSS_c_185_n N_ZI_c_271_n 4.67196e-19
cc_149 N_VSS_c_168_n N_ZI_c_276_n 2.68747e-19
cc_150 N_VSS_c_155_n N_ZI_c_277_n 3.44104e-19
cc_151 N_VSS_c_159_n N_ZI_c_277_n 5.20154e-19
cc_152 N_VSS_c_181_n N_ZI_c_277_n 8.7206e-19
cc_153 N_VSS_c_185_n N_ZI_c_277_n 0.0012589f
cc_154 N_VSS_c_179_n N_ZI_c_298_n 9.87505e-19
cc_155 N_VSS_c_148_n N_Z_c_329_n 3.43419e-19
cc_156 N_VSS_c_159_n N_Z_c_329_n 3.48267e-19
cc_157 N_VSS_c_148_n N_Z_c_332_n 3.48267e-19
cc_158 N_VSS_c_159_n N_Z_c_332_n 7.85754e-19
cc_159 N_VSS_c_227_p N_SELI_c_343_n 3.43419e-19
cc_160 N_VSS_c_150_n N_SELI_c_343_n 3.48267e-19
cc_161 N_VSS_c_227_p N_SELI_c_346_n 3.48267e-19
cc_162 N_VSS_c_150_n N_SELI_c_346_n 5.71987e-19
cc_163 N_VSS_c_163_n N_SELI_c_349_n 7.9573e-19
cc_164 N_VSS_c_175_n N_SELI_c_349_n 3.2351e-19
cc_165 N_VSS_c_188_n N_SELI_c_349_n 4.51137e-19
cc_166 N_VSS_c_194_n N_SELI_c_349_n 6.69121e-19
cc_167 N_VSS_c_159_n N_SELI_c_352_n 0.00105826f
cc_168 N_VSS_c_181_n N_SELI_c_352_n 3.89038e-19
cc_169 N_VSS_c_163_n N_SELI_c_368_n 3.2351e-19
cc_170 N_VSS_c_175_n N_SELI_c_368_n 0.00117301f
cc_171 N_VSS_c_188_n N_SELI_c_370_n 7.32115e-19
cc_172 N_VSS_c_194_n N_SELI_c_370_n 6.85767e-19
cc_173 N_VSS_XI7.X0_PGD N_SEL_c_419_n 3.9807e-19
cc_174 N_VSS_c_171_n N_SEL_c_430_n 9.4551e-19
cc_175 N_VSS_c_194_n N_SEL_c_421_n 2.60801e-19
cc_176 N_VSS_c_188_n N_SEL_c_422_n 2.64936e-19
cc_177 N_VSS_c_155_n N_SEL_c_433_n 3.36692e-19
cc_178 N_VSS_c_171_n N_SEL_c_433_n 3.29317e-19
cc_179 N_VSS_c_185_n N_SEL_c_425_n 3.72478e-19
cc_180 N_VSS_c_155_n N_SEL_c_427_n 3.2351e-19
cc_181 N_VSS_c_171_n N_SEL_c_427_n 2.68747e-19
cc_182 N_VSS_XI7.X0_PGS N_B_XI11.X0_PGS 0.00187616f
cc_183 N_VSS_XI9.X0_PGD N_B_XI11.X0_PGS 0.00145666f
cc_184 N_VSS_c_252_p N_B_c_495_n 0.00187616f
cc_185 N_VSS_c_163_n B 3.92469e-19
cc_186 N_VSS_c_175_n B 3.5189e-19
cc_187 N_VSS_c_185_n B 2.02689e-19
cc_188 N_VSS_XI9.X0_PGD N_B_c_491_n 3.23173e-19
cc_189 N_VSS_c_147_n N_B_c_491_n 0.00295829f
cc_190 N_VSS_c_163_n N_B_c_491_n 3.5189e-19
cc_191 N_VSS_c_171_n N_B_c_491_n 6.40394e-19
cc_192 N_VSS_c_175_n N_B_c_491_n 6.81736e-19
cc_193 N_VSS_c_188_n A 2.20363e-19
cc_194 N_ZI_c_262_n N_Z_c_329_n 6.8653e-19
cc_195 N_ZI_c_271_n N_SELI_c_346_n 6.18319e-19
cc_196 N_ZI_c_277_n N_SELI_c_346_n 0.00222064f
cc_197 N_ZI_c_262_n N_SELI_c_374_n 2.5026e-19
cc_198 N_ZI_c_283_n N_SELI_c_374_n 0.00194838f
cc_199 N_ZI_c_276_n N_SELI_c_374_n 9.76295e-19
cc_200 N_ZI_c_271_n N_SELI_c_349_n 0.00164769f
cc_201 N_ZI_c_269_n N_SELI_c_350_n 0.00166258f
cc_202 N_ZI_c_277_n N_SELI_c_350_n 0.00145462f
cc_203 N_ZI_c_262_n N_SELI_c_352_n 7.59552e-19
cc_204 N_ZI_c_277_n N_SELI_c_352_n 0.00172184f
cc_205 N_ZI_c_269_n N_SELI_c_370_n 7.67117e-19
cc_206 N_ZI_c_277_n N_SELI_c_370_n 7.85627e-19
cc_207 N_ZI_c_269_n N_SELI_c_384_n 6.01706e-19
cc_208 N_ZI_c_271_n N_SELI_c_384_n 3.05282e-19
cc_209 N_ZI_c_314_p N_SELI_c_384_n 6.45182e-19
cc_210 N_ZI_c_271_n N_SELI_c_387_n 8.23018e-19
cc_211 N_ZI_c_262_n N_SEL_c_419_n 0.00374573f
cc_212 N_ZI_c_276_n N_SEL_c_439_n 4.8006e-19
cc_213 N_ZI_c_264_n N_SEL_c_420_n 9.00465e-19
cc_214 N_ZI_c_271_n N_SEL_c_420_n 0.00250758f
cc_215 N_ZI_c_277_n N_SEL_c_420_n 8.4167e-19
cc_216 N_ZI_c_269_n N_SEL_c_421_n 9.51454e-19
cc_217 N_ZI_c_271_n N_SEL_c_421_n 4.59089e-19
cc_218 N_ZI_c_314_p N_SEL_c_421_n 0.00107464f
cc_219 N_ZI_c_263_n N_SEL_c_446_n 9.00465e-19
cc_220 N_ZI_c_269_n N_SEL_c_446_n 0.00242724f
cc_221 N_ZI_c_277_n N_SEL_c_433_n 0.0014877f
cc_222 N_ZI_c_262_n N_SEL_c_427_n 5.45742e-19
cc_223 N_ZI_XI4.X0_CG N_B_XI11.X0_PGS 0.00184555f
cc_224 N_Z_c_329_n N_SELI_c_374_n 7.7787e-19
cc_225 N_Z_c_332_n N_SELI_c_374_n 0.00121421f
cc_226 N_SELI_c_343_n N_SEL_c_419_n 6.8653e-19
cc_227 N_SELI_c_346_n N_SEL_c_419_n 8.57466e-19
cc_228 N_SELI_c_349_n N_SEL_c_420_n 0.00141479f
cc_229 N_SELI_c_368_n N_SEL_c_420_n 9.76295e-19
cc_230 N_SELI_c_346_n N_SEL_c_421_n 3.66824e-19
cc_231 N_SELI_c_350_n N_SEL_c_446_n 0.00170409f
cc_232 N_SELI_c_356_n N_SEL_c_446_n 9.29204e-19
cc_233 N_SELI_c_349_n N_SEL_c_422_n 9.45347e-19
cc_234 N_SELI_c_368_n N_SEL_c_422_n 4.56568e-19
cc_235 N_SELI_c_346_n N_SEL_c_433_n 0.00216212f
cc_236 N_SELI_c_352_n N_SEL_c_433_n 7.61973e-19
cc_237 N_SELI_c_352_n N_SEL_c_425_n 0.00193122f
cc_238 N_SELI_c_350_n N_SEL_c_462_n 0.00200661f
cc_239 N_SELI_c_346_n N_SEL_c_427_n 0.00109331f
cc_240 N_SELI_c_352_n N_SEL_c_427_n 4.73568e-19
cc_241 N_SELI_c_349_n N_SEL_c_465_n 3.48267e-19
cc_242 N_SELI_c_350_n N_SEL_c_465_n 4.95293e-19
cc_243 N_SELI_c_356_n N_SEL_c_465_n 0.00480115f
cc_244 N_SELI_c_368_n N_SEL_c_465_n 9.11855e-19
cc_245 N_SELI_c_349_n N_SEL_c_428_n 4.56568e-19
cc_246 N_SELI_c_350_n N_SEL_c_428_n 3.48267e-19
cc_247 N_SELI_c_356_n N_SEL_c_428_n 9.03632e-19
cc_248 N_SELI_c_368_n N_SEL_c_428_n 0.00244546f
cc_249 N_SELI_XI11.X0_CG N_B_XI11.X0_PGS 4.83278e-19
cc_250 N_SELI_c_346_n N_B_XI11.X0_PGS 2.54355e-19
cc_251 N_SELI_c_352_n N_B_XI11.X0_PGS 8.44835e-19
cc_252 N_SELI_c_356_n N_B_XI11.X0_PGS 0.00126314f
cc_253 N_SELI_c_417_p N_A_XI10.X0_PGS 5.12461e-19
cc_254 N_SELI_c_368_n N_A_XI10.X0_PGS 0.001089f
cc_255 N_SEL_c_473_p N_B_XI11.X0_PGS 2.07014e-19
cc_256 N_SEL_c_474_p N_B_XI11.X0_PGS 4.77845e-19
cc_257 N_SEL_c_425_n N_B_XI11.X0_PGS 7.3526e-19
cc_258 N_SEL_c_427_n N_B_XI11.X0_PGS 0.00100354f
cc_259 N_SEL_c_465_n N_B_XI11.X0_PGS 0.00142122f
cc_260 N_SEL_c_462_n B 4.4727e-19
cc_261 N_SEL_c_465_n B 3.2351e-19
cc_262 N_SEL_c_462_n N_B_c_491_n 3.29317e-19
cc_263 N_SEL_c_465_n N_B_c_491_n 0.00119577f
cc_264 N_SEL_XI10.X0_CG N_A_XI10.X0_PGS 4.99479e-19
cc_265 N_SEL_c_428_n N_A_XI10.X0_PGS 0.001089f
cc_266 N_SEL_c_484_p N_A_c_537_n 9.37683e-19
cc_267 N_SEL_c_422_n A 4.54408e-19
cc_268 N_SEL_c_428_n A 3.2351e-19
cc_269 N_SEL_c_422_n N_A_c_527_n 3.2351e-19
cc_270 N_SEL_c_428_n N_A_c_527_n 2.68747e-19
cc_271 N_B_XI11.X0_PGS N_A_XI10.X0_PGS 0.00134425f
*
.ends
*
*
.subckt MUX2_HPNW8 A B S0 Y VDD VSS
xgate (VDD VSS Y S0 B A) G4_MUX2_N2
.ends
*
* File: G3_MUXI2_N2.pex.netlist
* Created: Wed Mar  9 15:09:58 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MUXI2_N2_VSS 2 4 6 8 10 12 14 29 39 51 55 60 63 68 73 78 83 92 101
+ 110 111 117 123 129 131 136 138 140 141 144 145 146 Vss
c82 146 Vss 4.28045e-19
c83 145 Vss 3.62111e-19
c84 144 Vss 3.75522e-19
c85 141 Vss 0.00260366f
c86 138 Vss 0.00496506f
c87 136 Vss 0.00156482f
c88 131 Vss 0.00130885f
c89 129 Vss 0.0025874f
c90 124 Vss 0.00128107f
c91 123 Vss 0.00657991f
c92 117 Vss 0.0039834f
c93 111 Vss 0.00549375f
c94 110 Vss 0.0044599f
c95 101 Vss 0.00833837f
c96 92 Vss 0.0039597f
c97 83 Vss 2.73987e-19
c98 78 Vss 0.00101545f
c99 73 Vss 0.00217935f
c100 68 Vss 1.35342e-19
c101 63 Vss 7.10513e-22
c102 60 Vss 0.00389683f
c103 55 Vss 0.0017936f
c104 51 Vss 0.00537538f
c105 45 Vss 0.0783825f
c106 39 Vss 0.0354115f
c107 38 Vss 0.0688416f
c108 29 Vss 0.0347733f
c109 28 Vss 0.100982f
c110 14 Vss 0.135207f
c111 10 Vss 0.135463f
c112 6 Vss 0.135561f
c113 4 Vss 0.134971f
r114 137 146 0.551426
r115 137 138 15.5878
r116 136 146 0.551426
r117 135 136 4.58464
r118 131 146 0.0828784
r119 130 145 0.494161
r120 129 138 0.652036
r121 129 130 4.41793
r122 125 145 0.128424
r123 123 135 0.652036
r124 123 124 13.0037
r125 119 124 0.652036
r126 118 144 0.494161
r127 117 145 0.494161
r128 117 118 10.2946
r129 113 144 0.128424
r130 112 140 0.326018
r131 111 144 0.494161
r132 111 112 10.1279
r133 110 140 0.326018
r134 109 141 0.14525
r135 109 110 4.54296
r136 83 131 1.82344
r137 78 101 1.16709
r138 78 125 2.16729
r139 73 119 5.2515
r140 68 92 1.16709
r141 68 113 2.16729
r142 63 141 2.334
r143 60 83 1.16709
r144 55 73 1.16709
r145 51 63 1.16709
r146 45 101 0.0476429
r147 43 45 1.8672
r148 40 43 0.0685365
r149 38 43 0.5835
r150 38 39 2.8008
r151 35 39 0.652036
r152 31 92 0.0476429
r153 29 31 1.45875
r154 28 32 0.652036
r155 28 31 1.45875
r156 25 29 0.652036
r157 14 40 3.8511
r158 12 60 0.185659
r159 10 35 3.8511
r160 8 55 0.185659
r161 6 32 3.8511
r162 4 25 3.8511
r163 2 51 0.185659
.ends

.subckt PM_G3_MUXI2_N2_VDD 2 4 6 8 10 12 14 28 38 52 56 60 62 63 66 68 72 74 75
+ 76 80 81 83 84 86 87 89 98 Vss
c93 98 Vss 0.0111581f
c94 89 Vss 0.0046197f
c95 87 Vss 4.52364e-19
c96 84 Vss 4.42749e-19
c97 83 Vss 0.0021109f
c98 81 Vss 0.00811581f
c99 80 Vss 8.64091e-19
c100 76 Vss 0.00179444f
c101 75 Vss 6.09322e-19
c102 74 Vss 0.00543501f
c103 72 Vss 0.00102525f
c104 68 Vss 0.00843754f
c105 66 Vss 0.00123499f
c106 63 Vss 6.1175e-19
c107 62 Vss 0.00356077f
c108 60 Vss 6.73464e-19
c109 56 Vss 0.00425172f
c110 52 Vss 0.00654171f
c111 44 Vss 1.28925e-19
c112 39 Vss 0.0805856f
c113 38 Vss 0.103898f
c114 29 Vss 0.0367217f
c115 28 Vss 0.101295f
c116 12 Vss 0.134871f
c117 10 Vss 0.00143442f
c118 8 Vss 0.136499f
c119 4 Vss 0.136393f
c120 2 Vss 0.13497f
r121 82 87 0.551426
r122 82 83 4.58464
r123 81 87 0.551426
r124 80 86 0.326018
r125 80 81 15.5878
r126 76 87 0.0828784
r127 76 78 1.82344
r128 74 86 0.326018
r129 74 75 10.1279
r130 72 98 1.16709
r131 70 75 0.652036
r132 70 72 2.16729
r133 69 84 0.494161
r134 68 83 0.652036
r135 68 69 13.0037
r136 64 84 0.128424
r137 64 66 5.2515
r138 62 84 0.494161
r139 62 63 7.46046
r140 60 89 1.16709
r141 58 63 0.652036
r142 58 60 2.16729
r143 56 78 1.16709
r144 52 66 1.16709
r145 44 98 0.0476429
r146 44 46 1.92555
r147 39 46 0.5835
r148 38 40 0.652036
r149 38 39 2.8008
r150 35 46 0.0685365
r151 31 89 0.0476429
r152 29 31 1.45875
r153 28 32 0.652036
r154 28 31 1.45875
r155 25 29 0.652036
r156 14 56 0.185659
r157 12 40 3.8511
r158 10 52 0.185659
r159 8 35 3.8511
r160 6 52 0.185659
r161 4 25 3.8511
r162 2 32 3.8511
.ends

.subckt PM_G3_MUXI2_N2_SELI 2 4 6 8 21 29 33 35 38 43 53 58 72 77 78 Vss
c64 78 Vss 8.06863e-19
c65 72 Vss 0.00199393f
c66 58 Vss 0.00224258f
c67 53 Vss 0.00245485f
c68 43 Vss 9.25008e-19
c69 38 Vss 0.00141078f
c70 36 Vss 0.00169592f
c71 35 Vss 0.00419199f
c72 33 Vss 0.00348196f
c73 29 Vss 0.00522942f
c74 21 Vss 0.112066f
c75 6 Vss 0.112066f
c76 4 Vss 0.00143442f
r77 77 78 0.655813
r78 76 77 3.501
r79 72 76 0.655813
r80 43 53 1.16709
r81 43 72 2.00578
r82 43 46 0.333429
r83 38 58 1.16709
r84 38 78 2.00578
r85 35 46 0.0685365
r86 35 36 7.46046
r87 31 36 0.652036
r88 31 33 7.002
r89 29 33 1.16709
r90 21 58 0.50025
r91 18 53 0.50025
r92 8 21 3.09255
r93 6 18 3.09255
r94 4 29 0.185659
r95 2 29 0.185659
.ends

.subckt PM_G3_MUXI2_N2_SEL 2 4 6 8 16 22 26 37 40 42 46 51 58 63 68 72 77 78 Vss
c64 78 Vss 7.50288e-20
c65 77 Vss 9.69437e-20
c66 72 Vss 8.26714e-19
c67 68 Vss 0.00220099f
c68 63 Vss 0.00251571f
c69 58 Vss 0.00247916f
c70 51 Vss 3.96204e-19
c71 46 Vss 8.47469e-20
c72 42 Vss 0.00123172f
c73 37 Vss 0.00197358f
c74 26 Vss 0.11221f
c75 22 Vss 0.125771f
c76 20 Vss 0.0247918f
c77 17 Vss 0.036952f
c78 16 Vss 0.188224f
c79 8 Vss 0.112066f
c80 2 Vss 0.139232f
r81 76 78 0.655813
r82 76 77 3.501
r83 72 77 0.655813
r84 54 63 1.16709
r85 54 72 2.00578
r86 51 54 0.5835
r87 49 58 1.16709
r88 46 49 0.5835
r89 42 68 1.16709
r90 42 78 2.00578
r91 38 46 0.0685365
r92 38 40 1.45875
r93 37 51 0.0685365
r94 37 40 3.12589
r95 36 58 0.0476429
r96 33 68 0.50025
r97 26 63 0.50025
r98 22 58 0.357321
r99 20 36 0.326018
r100 20 22 0.40845
r101 17 36 6.7686
r102 16 36 0.326018
r103 16 36 0.1167
r104 13 17 0.652036
r105 8 33 3.09255
r106 6 26 3.09255
r107 4 22 3.44265
r108 2 13 3.8511
.ends

.subckt PM_G3_MUXI2_N2_B 2 4 7 16 20 24 27 Vss
c24 27 Vss 0.00705011f
c25 24 Vss 6.61761e-19
c26 20 Vss 0.0287936f
c27 16 Vss 0.0658163f
c28 7 Vss 0.142266f
c29 4 Vss 0.349678f
c30 2 Vss 0.11635f
r31 24 27 1.16709
r32 16 27 0.50025
r33 16 18 1.9839
r34 12 20 0.494161
r35 9 20 0.494161
r36 8 18 0.0685365
r37 7 20 0.128424
r38 7 8 4.7847
r39 4 12 11.0281
r40 2 9 3.20925
.ends

.subckt PM_G3_MUXI2_N2_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00368622f
c33 27 Vss 0.00747653f
c34 23 Vss 0.00756091f
c35 8 Vss 0.00143442f
c36 6 Vss 0.00143442f
r37 33 35 5.91836
r38 30 33 5.08479
r39 27 35 1.16709
r40 23 30 1.16709
r41 8 27 0.185659
r42 6 23 0.185659
r43 4 27 0.185659
r44 2 23 0.185659
.ends

.subckt PM_G3_MUXI2_N2_A 2 4 14 17 23 Vss
c23 23 Vss 0.00453252f
c24 17 Vss 3.94005e-19
c25 14 Vss 0.0840432f
c26 12 Vss 1.30835e-19
c27 2 Vss 0.557463f
r28 20 23 1.16709
r29 17 20 0.0416786
r30 12 23 0.0476429
r31 12 14 1.92555
r32 7 14 0.0685365
r33 2 4 15.4044
r34 2 7 3.8511
.ends

.subckt G3_MUXI2_N2  VSS VDD SEL B Z A
*
* A	A
* Z	Z
* B	B
* SEL	SEL
* VDD	VDD
* VSS	VSS
XI6.X0 N_SELI_XI6.X0_D N_VDD_XI6.X0_PGD N_SEL_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW8
XI7.X0 N_SELI_XI7.X0_D N_VSS_XI7.X0_PGD N_SEL_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW8
XI11.X0 N_Z_XI11.X0_D N_VDD_XI11.X0_PGD N_SELI_XI11.X0_CG N_B_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW8
XI9.X0 N_Z_XI9.X0_D N_VSS_XI9.X0_PGD N_SEL_XI9.X0_CG N_B_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW8
XI10.X0 N_Z_XI10.X0_D N_VDD_XI10.X0_PGD N_SEL_XI10.X0_CG N_A_XI10.X0_PGS
+ N_VSS_XI10.X0_S TIGFET_HPNW8
XI8.X0 N_Z_XI8.X0_D N_VSS_XI8.X0_PGD N_SELI_XI8.X0_CG N_A_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW8
*
x_PM_G3_MUXI2_N2_VSS N_VSS_XI6.X0_S N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS
+ N_VSS_XI11.X0_S N_VSS_XI9.X0_PGD N_VSS_XI10.X0_S N_VSS_XI8.X0_PGD N_VSS_c_4_p
+ N_VSS_c_20_p N_VSS_c_45_p N_VSS_c_72_p N_VSS_c_27_p N_VSS_c_46_p N_VSS_c_5_p
+ N_VSS_c_26_p N_VSS_c_17_p N_VSS_c_28_p N_VSS_c_9_p N_VSS_c_19_p N_VSS_c_6_p
+ N_VSS_c_10_p N_VSS_c_11_p N_VSS_c_29_p N_VSS_c_24_p N_VSS_c_31_p N_VSS_c_34_p
+ N_VSS_c_35_p VSS N_VSS_c_50_p N_VSS_c_12_p N_VSS_c_25_p N_VSS_c_36_p Vss
+ PM_G3_MUXI2_N2_VSS
x_PM_G3_MUXI2_N2_VDD N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI7.X0_S
+ N_VDD_XI11.X0_PGD N_VDD_XI9.X0_S N_VDD_XI10.X0_PGD N_VDD_XI8.X0_S N_VDD_c_86_n
+ N_VDD_c_171_p N_VDD_c_127_p N_VDD_c_151_p N_VDD_c_87_n N_VDD_c_89_n
+ N_VDD_c_95_n N_VDD_c_96_n N_VDD_c_102_n N_VDD_c_108_n N_VDD_c_109_n
+ N_VDD_c_112_n N_VDD_c_113_n N_VDD_c_114_n N_VDD_c_115_n N_VDD_c_119_n
+ N_VDD_c_122_n VDD N_VDD_c_123_n N_VDD_c_124_n N_VDD_c_126_n Vss
+ PM_G3_MUXI2_N2_VDD
x_PM_G3_MUXI2_N2_SELI N_SELI_XI6.X0_D N_SELI_XI7.X0_D N_SELI_XI11.X0_CG
+ N_SELI_XI8.X0_CG N_SELI_c_238_p N_SELI_c_176_n N_SELI_c_178_n N_SELI_c_182_n
+ N_SELI_c_183_n N_SELI_c_197_n N_SELI_c_199_n N_SELI_c_186_n N_SELI_c_188_n
+ N_SELI_c_189_n N_SELI_c_220_p Vss PM_G3_MUXI2_N2_SELI
x_PM_G3_MUXI2_N2_SEL N_SEL_XI6.X0_CG N_SEL_XI7.X0_CG N_SEL_XI9.X0_CG
+ N_SEL_XI10.X0_CG N_SEL_c_240_n N_SEL_c_283_p N_SEL_c_284_p N_SEL_c_241_n SEL
+ N_SEL_c_242_n N_SEL_c_243_n N_SEL_c_256_n N_SEL_c_245_n N_SEL_c_271_n
+ N_SEL_c_257_n N_SEL_c_247_n N_SEL_c_249_n N_SEL_c_250_n Vss PM_G3_MUXI2_N2_SEL
x_PM_G3_MUXI2_N2_B N_B_XI11.X0_PGS N_B_XI9.X0_PGS N_B_c_304_n N_B_c_324_n
+ N_B_c_315_n B N_B_c_306_n Vss PM_G3_MUXI2_N2_B
x_PM_G3_MUXI2_N2_Z N_Z_XI11.X0_D N_Z_XI9.X0_D N_Z_XI10.X0_D N_Z_XI8.X0_D
+ N_Z_c_328_n N_Z_c_338_n N_Z_c_332_n Z Vss PM_G3_MUXI2_N2_Z
x_PM_G3_MUXI2_N2_A N_A_XI10.X0_PGS N_A_XI8.X0_PGS N_A_c_362_n A N_A_c_368_n Vss
+ PM_G3_MUXI2_N2_A
cc_1 N_VSS_XI7.X0_PGD N_VDD_XI6.X0_PGD 0.00200584f
cc_2 N_VSS_XI9.X0_PGD N_VDD_XI11.X0_PGD 2.37403e-19
cc_3 N_VSS_XI8.X0_PGD N_VDD_XI10.X0_PGD 2.37403e-19
cc_4 N_VSS_c_4_p N_VDD_c_86_n 0.00200584f
cc_5 N_VSS_c_5_p N_VDD_c_87_n 7.57561e-19
cc_6 N_VSS_c_6_p N_VDD_c_87_n 8.35657e-19
cc_7 N_VSS_c_4_p N_VDD_c_89_n 3.9313e-19
cc_8 N_VSS_c_5_p N_VDD_c_89_n 0.00161703f
cc_9 N_VSS_c_9_p N_VDD_c_89_n 2.26455e-19
cc_10 N_VSS_c_10_p N_VDD_c_89_n 0.0043279f
cc_11 N_VSS_c_11_p N_VDD_c_89_n 0.00126887f
cc_12 N_VSS_c_12_p N_VDD_c_89_n 7.74609e-19
cc_13 N_VSS_c_10_p N_VDD_c_95_n 0.00157719f
cc_14 N_VSS_XI7.X0_PGS N_VDD_c_96_n 2.59535e-19
cc_15 N_VSS_XI9.X0_PGD N_VDD_c_96_n 2.19376e-19
cc_16 N_VSS_c_5_p N_VDD_c_96_n 0.00180638f
cc_17 N_VSS_c_17_p N_VDD_c_96_n 7.4365e-19
cc_18 N_VSS_c_9_p N_VDD_c_96_n 9.55109e-19
cc_19 N_VSS_c_19_p N_VDD_c_96_n 2.70301e-19
cc_20 N_VSS_c_20_p N_VDD_c_102_n 0.00111089f
cc_21 N_VSS_c_17_p N_VDD_c_102_n 0.00161703f
cc_22 N_VSS_c_19_p N_VDD_c_102_n 2.26455e-19
cc_23 N_VSS_c_11_p N_VDD_c_102_n 0.00574413f
cc_24 N_VSS_c_24_p N_VDD_c_102_n 0.00456934f
cc_25 N_VSS_c_25_p N_VDD_c_102_n 7.61747e-19
cc_26 N_VSS_c_26_p N_VDD_c_108_n 0.00121523f
cc_27 N_VSS_c_27_p N_VDD_c_109_n 3.4118e-19
cc_28 N_VSS_c_28_p N_VDD_c_109_n 4.19648e-19
cc_29 N_VSS_c_29_p N_VDD_c_109_n 0.00755466f
cc_30 N_VSS_c_29_p N_VDD_c_112_n 0.00152669f
cc_31 N_VSS_c_31_p N_VDD_c_113_n 4.68065e-19
cc_32 N_VSS_c_29_p N_VDD_c_114_n 0.00106538f
cc_33 N_VSS_c_28_p N_VDD_c_115_n 0.00187494f
cc_34 N_VSS_c_34_p N_VDD_c_115_n 0.00339451f
cc_35 N_VSS_c_35_p N_VDD_c_115_n 0.00671233f
cc_36 N_VSS_c_36_p N_VDD_c_115_n 9.16632e-19
cc_37 N_VSS_c_17_p N_VDD_c_119_n 4.28751e-19
cc_38 N_VSS_c_19_p N_VDD_c_119_n 3.63088e-19
cc_39 N_VSS_c_35_p N_VDD_c_119_n 0.00337584f
cc_40 N_VSS_c_11_p N_VDD_c_122_n 0.0011585f
cc_41 N_VSS_c_35_p N_VDD_c_123_n 0.00100712f
cc_42 N_VSS_c_5_p N_VDD_c_124_n 3.48267e-19
cc_43 N_VSS_c_9_p N_VDD_c_124_n 6.46219e-19
cc_44 N_VSS_c_26_p N_VDD_c_126_n 2.84469e-19
cc_45 N_VSS_c_45_p N_SELI_c_176_n 3.43419e-19
cc_46 N_VSS_c_46_p N_SELI_c_176_n 3.48267e-19
cc_47 N_VSS_c_45_p N_SELI_c_178_n 3.48267e-19
cc_48 N_VSS_c_46_p N_SELI_c_178_n 5.71987e-19
cc_49 N_VSS_c_10_p N_SELI_c_178_n 2.50156e-19
cc_50 N_VSS_c_50_p N_SELI_c_178_n 2.7826e-19
cc_51 N_VSS_c_26_p N_SELI_c_182_n 0.00111908f
cc_52 N_VSS_c_17_p N_SELI_c_183_n 8.64455e-19
cc_53 N_VSS_c_19_p N_SELI_c_183_n 3.49905e-19
cc_54 N_VSS_c_35_p N_SELI_c_183_n 9.07743e-19
cc_55 N_VSS_c_17_p N_SELI_c_186_n 3.2351e-19
cc_56 N_VSS_c_19_p N_SELI_c_186_n 2.68747e-19
cc_57 N_VSS_c_29_p N_SELI_c_188_n 6.74415e-19
cc_58 N_VSS_c_35_p N_SELI_c_189_n 5.03655e-19
cc_59 N_VSS_XI7.X0_PGD N_SEL_c_240_n 4.18141e-19
cc_60 N_VSS_c_11_p N_SEL_c_241_n 5.08457e-19
cc_61 N_VSS_c_35_p N_SEL_c_242_n 7.91494e-19
cc_62 N_VSS_c_5_p N_SEL_c_243_n 5.97048e-19
cc_63 N_VSS_c_9_p N_SEL_c_243_n 3.08902e-19
cc_64 N_VSS_c_5_p N_SEL_c_245_n 3.2351e-19
cc_65 N_VSS_c_9_p N_SEL_c_245_n 2.68747e-19
cc_66 N_VSS_c_11_p N_SEL_c_247_n 0.00100236f
cc_67 N_VSS_c_29_p N_SEL_c_247_n 2.48958e-19
cc_68 N_VSS_c_35_p N_SEL_c_249_n 4.36463e-19
cc_69 N_VSS_c_29_p N_SEL_c_250_n 9.32613e-19
cc_70 N_VSS_XI7.X0_PGS N_B_c_304_n 2.56596e-19
cc_71 N_VSS_c_26_p B 0.00157463f
cc_72 N_VSS_c_72_p N_B_c_306_n 0.00246958f
cc_73 N_VSS_c_26_p N_B_c_306_n 8.835e-19
cc_74 N_VSS_c_72_p N_Z_c_328_n 3.43419e-19
cc_75 N_VSS_c_27_p N_Z_c_328_n 3.43419e-19
cc_76 N_VSS_c_26_p N_Z_c_328_n 3.48267e-19
cc_77 N_VSS_c_28_p N_Z_c_328_n 3.48267e-19
cc_78 N_VSS_c_72_p N_Z_c_332_n 3.48267e-19
cc_79 N_VSS_c_27_p N_Z_c_332_n 3.48267e-19
cc_80 N_VSS_c_26_p N_Z_c_332_n 5.71987e-19
cc_81 N_VSS_c_28_p N_Z_c_332_n 5.71987e-19
cc_82 N_VSS_c_35_p N_Z_c_332_n 6.72116e-19
cc_83 N_VDD_c_127_p N_SELI_c_176_n 3.43419e-19
cc_84 N_VDD_c_89_n N_SELI_c_176_n 3.4118e-19
cc_85 N_VDD_c_96_n N_SELI_c_176_n 3.48267e-19
cc_86 N_VDD_c_127_p N_SELI_c_178_n 3.48267e-19
cc_87 N_VDD_c_89_n N_SELI_c_178_n 4.78806e-19
cc_88 N_VDD_c_96_n N_SELI_c_178_n 7.09569e-19
cc_89 N_VDD_c_115_n N_SELI_c_183_n 6.15494e-19
cc_90 N_VDD_c_108_n N_SELI_c_197_n 4.44319e-19
cc_91 N_VDD_c_126_n N_SELI_c_197_n 3.49905e-19
cc_92 N_VDD_c_108_n N_SELI_c_199_n 3.43988e-19
cc_93 N_VDD_c_126_n N_SELI_c_199_n 2.68747e-19
cc_94 N_VDD_c_115_n N_SELI_c_186_n 3.66936e-19
cc_95 N_VDD_XI6.X0_PGD N_SEL_c_240_n 4.28909e-19
cc_96 N_VDD_c_127_p N_SEL_c_241_n 6.34806e-19
cc_97 N_VDD_c_96_n N_SEL_c_241_n 0.00105602f
cc_98 N_VDD_c_109_n N_SEL_c_242_n 2.67421e-19
cc_99 N_VDD_c_115_n N_SEL_c_242_n 6.15494e-19
cc_100 N_VDD_c_102_n N_SEL_c_256_n 2.25302e-19
cc_101 N_VDD_c_115_n N_SEL_c_257_n 3.66936e-19
cc_102 N_VDD_c_102_n N_SEL_c_247_n 4.27423e-19
cc_103 N_VDD_c_115_n N_SEL_c_249_n 2.2501e-19
cc_104 N_VDD_c_127_p N_B_c_304_n 2.2574e-19
cc_105 N_VDD_c_109_n N_Z_c_328_n 3.4118e-19
cc_106 N_VDD_c_127_p N_Z_c_338_n 3.43419e-19
cc_107 N_VDD_c_151_p N_Z_c_338_n 3.43419e-19
cc_108 N_VDD_c_96_n N_Z_c_338_n 3.48267e-19
cc_109 N_VDD_c_102_n N_Z_c_338_n 3.4118e-19
cc_110 N_VDD_c_113_n N_Z_c_338_n 3.72199e-19
cc_111 N_VDD_c_127_p N_Z_c_332_n 3.48267e-19
cc_112 N_VDD_c_151_p N_Z_c_332_n 3.48267e-19
cc_113 N_VDD_c_96_n N_Z_c_332_n 8.16241e-19
cc_114 N_VDD_c_102_n N_Z_c_332_n 4.7984e-19
cc_115 N_VDD_c_109_n N_Z_c_332_n 4.7984e-19
cc_116 N_VDD_c_113_n N_Z_c_332_n 8.08807e-19
cc_117 N_VDD_c_115_n N_Z_c_332_n 9.6188e-19
cc_118 N_VDD_XI10.X0_PGD N_A_XI10.X0_PGS 0.00151037f
cc_119 N_VDD_c_115_n N_A_XI10.X0_PGS 0.00102341f
cc_120 N_VDD_c_109_n N_A_c_362_n 3.60536e-19
cc_121 N_VDD_c_115_n N_A_c_362_n 3.92733e-19
cc_122 N_VDD_c_108_n A 5.33592e-19
cc_123 N_VDD_c_109_n A 0.00141439f
cc_124 N_VDD_c_115_n A 5.00176e-19
cc_125 N_VDD_c_126_n A 3.48267e-19
cc_126 N_VDD_XI10.X0_PGD N_A_c_368_n 3.23173e-19
cc_127 N_VDD_c_171_p N_A_c_368_n 0.00480616f
cc_128 N_VDD_c_108_n N_A_c_368_n 4.04186e-19
cc_129 N_VDD_c_109_n N_A_c_368_n 0.00120343f
cc_130 N_VDD_c_115_n N_A_c_368_n 3.66936e-19
cc_131 N_VDD_c_126_n N_A_c_368_n 6.39485e-19
cc_132 N_SELI_c_176_n N_SEL_c_240_n 6.55689e-19
cc_133 N_SELI_c_178_n N_SEL_c_240_n 9.27181e-19
cc_134 N_SELI_c_182_n N_SEL_c_240_n 4.08878e-19
cc_135 N_SELI_c_197_n N_SEL_c_241_n 0.00289751f
cc_136 N_SELI_c_183_n N_SEL_c_242_n 0.00240159f
cc_137 N_SELI_c_186_n N_SEL_c_242_n 4.99367e-19
cc_138 N_SELI_c_178_n N_SEL_c_243_n 0.0024269f
cc_139 N_SELI_c_182_n N_SEL_c_243_n 0.00289751f
cc_140 N_SELI_c_199_n N_SEL_c_256_n 5.42085e-19
cc_141 N_SELI_c_178_n N_SEL_c_245_n 0.00100994f
cc_142 N_SELI_c_182_n N_SEL_c_245_n 5.66159e-19
cc_143 N_SELI_c_199_n N_SEL_c_271_n 0.00493717f
cc_144 N_SELI_c_186_n N_SEL_c_271_n 8.7809e-19
cc_145 N_SELI_c_199_n N_SEL_c_257_n 8.69867e-19
cc_146 N_SELI_c_186_n N_SEL_c_257_n 0.00494248f
cc_147 N_SELI_c_183_n N_SEL_c_247_n 0.00165721f
cc_148 N_SELI_c_197_n N_SEL_c_247_n 4.7869e-19
cc_149 N_SELI_c_188_n N_SEL_c_247_n 9.53674e-19
cc_150 N_SELI_c_220_p N_SEL_c_247_n 7.98252e-19
cc_151 N_SELI_c_178_n N_SEL_c_249_n 3.01017e-19
cc_152 N_SELI_c_189_n N_SEL_c_249_n 0.00144491f
cc_153 N_SELI_c_197_n N_SEL_c_250_n 0.00165436f
cc_154 N_SELI_c_188_n N_SEL_c_250_n 7.97695e-19
cc_155 N_SELI_XI11.X0_CG N_B_XI11.X0_PGS 4.31731e-19
cc_156 N_SELI_c_199_n N_B_XI11.X0_PGS 6.66106e-19
cc_157 N_SELI_c_178_n N_B_XI9.X0_PGS 2.97793e-19
cc_158 N_SELI_c_182_n N_B_XI9.X0_PGS 3.99745e-19
cc_159 N_SELI_c_199_n N_B_XI9.X0_PGS 5.45575e-19
cc_160 N_SELI_c_182_n N_B_c_304_n 4.011e-19
cc_161 N_SELI_c_182_n N_B_c_315_n 5.40503e-19
cc_162 N_SELI_c_199_n N_B_c_315_n 0.00179467f
cc_163 N_SELI_c_182_n B 0.00128002f
cc_164 N_SELI_c_182_n N_B_c_306_n 0.00106912f
cc_165 N_SELI_c_178_n N_Z_c_332_n 8.31671e-19
cc_166 N_SELI_c_183_n N_Z_c_332_n 0.00208341f
cc_167 N_SELI_c_197_n N_Z_c_332_n 0.00213869f
cc_168 N_SELI_c_238_p N_A_XI10.X0_PGS 5.00154e-19
cc_169 N_SELI_c_186_n N_A_XI10.X0_PGS 0.00276355f
cc_170 N_SEL_c_283_p N_B_XI9.X0_PGS 2.04953e-19
cc_171 N_SEL_c_284_p N_B_XI9.X0_PGS 4.65537e-19
cc_172 N_SEL_c_241_n N_B_XI9.X0_PGS 8.3216e-19
cc_173 N_SEL_c_245_n N_B_XI9.X0_PGS 0.00100354f
cc_174 N_SEL_c_271_n N_B_XI9.X0_PGS 0.00202689f
cc_175 N_SEL_c_241_n N_B_c_324_n 2.88938e-19
cc_176 N_SEL_c_245_n N_B_c_324_n 7.65159e-19
cc_177 N_SEL_c_245_n N_B_c_306_n 8.68391e-19
cc_178 N_SEL_c_242_n N_Z_c_332_n 0.00189968f
cc_179 N_SEL_c_256_n N_Z_c_332_n 0.00221938f
cc_180 N_SEL_c_271_n N_Z_c_332_n 9.50991e-19
cc_181 N_SEL_c_257_n N_Z_c_332_n 9.35582e-19
cc_182 N_SEL_c_247_n N_Z_c_332_n 9.18344e-19
cc_183 N_SEL_c_249_n N_Z_c_332_n 0.0021646f
cc_184 N_SEL_c_250_n N_Z_c_332_n 9.04233e-19
cc_185 N_SEL_XI10.X0_CG N_A_XI10.X0_PGS 4.87172e-19
cc_186 N_SEL_c_257_n N_A_XI10.X0_PGS 0.00276355f
cc_187 N_SEL_c_242_n A 4.55825e-19
cc_188 N_SEL_c_257_n A 3.2351e-19
cc_189 N_SEL_c_242_n N_A_c_368_n 3.49905e-19
cc_190 N_SEL_c_257_n N_A_c_368_n 2.68747e-19
cc_191 N_B_XI11.X0_PGS N_A_XI10.X0_PGS 0.00134199f
*
.ends
*
*
.subckt MUXI2_HPNW8 A B S0 Y VDD VSS
xgate (VSS VDD S0 B Y A) G3_MUXI2_N2
.ends
*
* File: G2_NAND2_N2.pex.netlist
* Created: Fri Feb 25 16:38:49 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NAND2_N2_VSS 2 3 5 6 8 18 19 21 41 47 52 61 68 73 74 Vss
c28 74 Vss 8.01054e-19
c29 73 Vss 0.00222032f
c30 69 Vss 0.00133128f
c31 68 Vss 0.00979385f
c32 61 Vss 0.00460027f
c33 52 Vss 0.00163484f
c34 47 Vss 0.00135376f
c35 41 Vss 0.00500207f
c36 38 Vss 0.0299355f
c37 37 Vss 0.0299355f
c38 32 Vss 0.105904f
c39 26 Vss 0.0688517f
c40 21 Vss 5.38535e-20
c41 19 Vss 0.0340588f
c42 18 Vss 0.064644f
c43 8 Vss 0.138428f
c44 6 Vss 0.137392f
c45 5 Vss 0.138084f
c46 3 Vss 0.137146f
r47 73 75 0.652036
r48 73 74 4.33457
r49 66 74 0.652036
r50 66 68 7.66886
r51 65 69 0.655813
r52 65 68 8.96089
r53 52 61 1.16709
r54 52 75 2.16729
r55 47 69 1.82344
r56 41 47 1.16709
r57 33 38 0.494161
r58 32 34 0.652036
r59 32 33 2.9175
r60 28 38 0.128424
r61 27 37 0.494161
r62 26 38 0.494161
r63 26 27 2.8008
r64 22 37 0.128424
r65 21 61 0.238214
r66 19 21 1.4004
r67 18 37 0.494161
r68 18 21 1.5171
r69 15 19 0.652036
r70 8 34 3.8511
r71 6 28 3.8511
r72 5 15 3.8511
r73 3 22 3.8511
r74 2 41 0.185659
.ends

.subckt PM_G2_NAND2_N2_VDD 1 3 5 15 17 22 27 31 32 34 36 37 38 42 47 49 52 58
+ Vss
c41 58 Vss 0.00548438f
c42 50 Vss 9.22237e-19
c43 49 Vss 0.00628406f
c44 47 Vss 0.00776909f
c45 42 Vss 0.00125451f
c46 38 Vss 0.00692242f
c47 37 Vss 8.60438e-19
c48 36 Vss 0.0123084f
c49 34 Vss 0.00177187f
c50 32 Vss 8.19549e-19
c51 31 Vss 0.00243037f
c52 27 Vss 0.00484855f
c53 22 Vss 0.00385756f
c54 17 Vss 0.171989f
c55 15 Vss 0.0339269f
c56 1 Vss 0.117266f
r57 49 52 0.326018
r58 48 50 0.551426
r59 48 49 5.08479
r60 47 50 0.551426
r61 46 47 8.54411
r62 42 50 0.0828784
r63 42 44 1.82344
r64 40 58 1.16709
r65 38 46 0.655813
r66 38 40 4.37625
r67 36 52 0.326018
r68 36 37 15.6711
r69 32 34 1.76818
r70 31 37 0.652036
r71 30 32 0.657751
r72 30 31 5.04311
r73 27 44 1.16709
r74 22 34 1.16709
r75 17 58 0.428786
r76 15 17 5.3682
r77 11 15 0.652036
r78 5 27 0.185659
r79 3 22 0.185659
r80 1 11 3.1509
.ends

.subckt PM_G2_NAND2_N2_A 2 4 13 18 21 26 31 Vss
c20 31 Vss 0.00388303f
c21 26 Vss 0.00333046f
c22 18 Vss 0.00166538f
c23 13 Vss 0.112394f
c24 2 Vss 0.111896f
r25 23 31 1.16709
r26 21 23 2.54239
r27 18 26 1.16709
r28 18 21 2.83414
r29 13 31 0.50025
r30 10 26 0.50025
r31 4 13 3.09255
r32 2 10 3.09255
.ends

.subckt PM_G2_NAND2_N2_Z 2 4 6 18 22 25 28 Vss
c26 25 Vss 0.00212593f
c27 22 Vss 0.00585482f
c28 18 Vss 0.00354571f
c29 6 Vss 0.00143442f
r30 28 30 4.83471
r31 25 28 6.71025
r32 22 30 1.16709
r33 18 25 1.16709
r34 6 22 0.185659
r35 4 22 0.185659
r36 2 18 0.185659
.ends

.subckt PM_G2_NAND2_N2_B 2 4 10 11 14 18 21 Vss
c23 18 Vss 9.58314e-20
c24 14 Vss 0.181262f
c25 11 Vss 0.0357204f
c26 10 Vss 0.288966f
c27 2 Vss 0.281263f
r28 18 21 0.0416786
r29 14 18 1.16709
r30 12 14 2.1006
r31 10 12 0.652036
r32 10 11 8.92755
r33 7 11 0.652036
r34 4 14 4.3179
r35 2 7 8.57745
.ends

.subckt G2_NAND2_N2  VSS VDD A Z B
*
* B	B
* Z	Z
* A	A
* VDD	VDD
* VSS	VSS
XI12.X0 N_Z_XI12.X0_D N_VDD_XI12.X0_PGD N_A_XI12.X0_CG N_B_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW8
XI10.X0 N_Z_XI10.X0_D N_VSS_XI10.X0_PGD N_A_XI10.X0_CG N_VSS_XI10.X0_PGS
+ N_VDD_XI10.X0_S TIGFET_HPNW8
XI11.X0 N_Z_XI11.X0_D N_VSS_XI11.X0_PGD N_B_XI11.X0_CG N_VSS_XI11.X0_PGS
+ N_VDD_XI11.X0_S TIGFET_HPNW8
*
x_PM_G2_NAND2_N2_VSS N_VSS_XI12.X0_S N_VSS_XI10.X0_PGD N_VSS_XI10.X0_PGS
+ N_VSS_XI11.X0_PGD N_VSS_XI11.X0_PGS N_VSS_c_7_p N_VSS_c_8_p N_VSS_c_19_p
+ N_VSS_c_22_p N_VSS_c_6_p N_VSS_c_2_p N_VSS_c_3_p VSS N_VSS_c_11_p N_VSS_c_12_p
+ Vss PM_G2_NAND2_N2_VSS
x_PM_G2_NAND2_N2_VDD N_VDD_XI12.X0_PGD N_VDD_XI10.X0_S N_VDD_XI11.X0_S
+ N_VDD_c_62_p N_VDD_c_52_p N_VDD_c_47_p N_VDD_c_48_p N_VDD_c_29_n N_VDD_c_33_n
+ N_VDD_c_34_n N_VDD_c_35_n N_VDD_c_40_n N_VDD_c_57_p N_VDD_c_51_p N_VDD_c_59_p
+ N_VDD_c_41_n VDD N_VDD_c_45_p Vss PM_G2_NAND2_N2_VDD
x_PM_G2_NAND2_N2_A N_A_XI12.X0_CG N_A_XI10.X0_CG N_A_c_70_n N_A_c_71_n A
+ N_A_c_78_n N_A_c_74_n Vss PM_G2_NAND2_N2_A
x_PM_G2_NAND2_N2_Z N_Z_XI12.X0_D N_Z_XI10.X0_D N_Z_XI11.X0_D N_Z_c_90_n
+ N_Z_c_95_n N_Z_c_92_n Z Vss PM_G2_NAND2_N2_Z
x_PM_G2_NAND2_N2_B N_B_XI12.X0_PGS N_B_XI11.X0_CG N_B_c_116_n N_B_c_118_n
+ N_B_c_121_n N_B_c_124_n B Vss PM_G2_NAND2_N2_B
cc_1 N_VSS_XI10.X0_PGS N_VDD_c_29_n 2.7398e-19
cc_2 N_VSS_c_2_p N_VDD_c_29_n 4.50283e-19
cc_3 N_VSS_c_3_p N_VDD_c_29_n 3.70842e-19
cc_4 VSS N_VDD_c_29_n 0.00384148f
cc_5 VSS N_VDD_c_33_n 0.0016639f
cc_6 N_VSS_c_6_p N_VDD_c_34_n 4.48301e-19
cc_7 N_VSS_c_7_p N_VDD_c_35_n 0.00183557f
cc_8 N_VSS_c_8_p N_VDD_c_35_n 3.51214e-19
cc_9 N_VSS_c_2_p N_VDD_c_35_n 0.00161703f
cc_10 N_VSS_c_3_p N_VDD_c_35_n 2.03837e-19
cc_11 N_VSS_c_11_p N_VDD_c_35_n 0.00517826f
cc_12 N_VSS_c_12_p N_VDD_c_40_n 0.00104633f
cc_13 N_VSS_XI11.X0_PGS N_VDD_c_41_n 3.32059e-19
cc_14 N_VSS_c_2_p N_VDD_c_41_n 2.24202e-19
cc_15 N_VSS_c_3_p N_A_c_70_n 0.00249847f
cc_16 N_VSS_c_2_p N_A_c_71_n 2.94885e-19
cc_17 N_VSS_c_3_p N_A_c_71_n 3.71222e-19
cc_18 VSS N_A_c_71_n 0.00255481f
cc_19 N_VSS_c_19_p N_A_c_74_n 3.96531e-19
cc_20 N_VSS_c_2_p N_A_c_74_n 2.87758e-19
cc_21 N_VSS_c_3_p N_A_c_74_n 8.98435e-19
cc_22 N_VSS_c_22_p N_Z_c_90_n 3.43419e-19
cc_23 N_VSS_c_6_p N_Z_c_90_n 3.48267e-19
cc_24 N_VSS_c_6_p N_Z_c_92_n 8.92744e-19
cc_25 VSS N_Z_c_92_n 7.39325e-19
cc_26 N_VSS_XI10.X0_PGD N_B_c_116_n 8.28117e-19
cc_27 N_VSS_XI11.X0_PGD N_B_c_116_n 8.28117e-19
cc_28 N_VSS_XI10.X0_PGS N_B_c_118_n 9.94582e-19
cc_29 N_VDD_XI12.X0_PGD N_A_XI12.X0_CG 5.34714e-19
cc_30 N_VDD_XI12.X0_PGD N_A_c_78_n 2.78309e-19
cc_31 N_VDD_c_45_p N_A_c_78_n 4.44265e-19
cc_32 N_VDD_c_45_p N_Z_c_90_n 0.00132057f
cc_33 N_VDD_c_47_p N_Z_c_95_n 3.43419e-19
cc_34 N_VDD_c_48_p N_Z_c_95_n 3.43419e-19
cc_35 N_VDD_c_34_n N_Z_c_95_n 3.72199e-19
cc_36 N_VDD_c_35_n N_Z_c_95_n 3.02646e-19
cc_37 N_VDD_c_51_p N_Z_c_95_n 3.72199e-19
cc_38 N_VDD_c_52_p N_Z_c_92_n 8.40856e-19
cc_39 N_VDD_c_47_p N_Z_c_92_n 3.48267e-19
cc_40 N_VDD_c_48_p N_Z_c_92_n 3.48267e-19
cc_41 N_VDD_c_34_n N_Z_c_92_n 8.08807e-19
cc_42 N_VDD_c_35_n N_Z_c_92_n 5.981e-19
cc_43 N_VDD_c_57_p N_Z_c_92_n 0.00172841f
cc_44 N_VDD_c_51_p N_Z_c_92_n 8.49942e-19
cc_45 N_VDD_c_59_p N_Z_c_92_n 0.00179028f
cc_46 N_VDD_c_45_p N_Z_c_92_n 8.835e-19
cc_47 N_VDD_XI12.X0_PGD N_B_XI12.X0_PGS 0.00153438f
cc_48 N_VDD_c_62_p N_B_c_116_n 0.00429636f
cc_49 N_VDD_c_57_p N_B_c_121_n 2.79672e-19
cc_50 N_VDD_c_59_p N_B_c_121_n 5.52596e-19
cc_51 N_VDD_c_45_p N_B_c_121_n 7.42072e-19
cc_52 N_VDD_c_35_n N_B_c_124_n 3.13539e-19
cc_53 N_VDD_c_57_p N_B_c_124_n 3.88313e-19
cc_54 N_VDD_c_59_p N_B_c_124_n 6.60945e-19
cc_55 N_VDD_c_45_p N_B_c_124_n 2.79672e-19
cc_56 N_A_c_71_n N_Z_c_92_n 0.0082161f
cc_57 N_A_c_78_n N_Z_c_92_n 9.58524e-19
cc_58 N_A_c_74_n N_Z_c_92_n 0.00100714f
cc_59 N_A_XI12.X0_CG N_B_XI12.X0_PGS 5.00154e-19
cc_60 N_A_c_71_n N_B_XI12.X0_PGS 7.2582e-19
cc_61 N_A_c_78_n N_B_XI12.X0_PGS 5.6636e-19
cc_62 N_A_c_71_n N_B_c_116_n 3.15161e-19
cc_63 N_A_c_78_n N_B_c_116_n 7.2846e-19
cc_64 N_A_c_74_n N_B_c_116_n 0.00228839f
cc_65 N_A_c_74_n N_B_c_121_n 9.27569e-19
cc_66 N_Z_c_95_n N_B_c_116_n 3.74089e-19
cc_67 N_Z_c_92_n N_B_c_116_n 4.8079e-19
cc_68 N_Z_c_92_n N_B_c_121_n 0.00105292f
cc_69 N_Z_c_92_n N_B_c_124_n 0.00147455f
*
.ends
*
*
.subckt NAND2_HPNW8 A B Y VDD VSS
xgate (VSS VDD A Y B) G2_NAND2_N2
.ends
*
* File: G2_NOR2_N2.pex.netlist
* Created: Mon Feb 28 09:43:23 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NOR2_N2_VSS 2 4 6 18 23 28 31 36 41 50 59 60 64 65 70 77 78 80 Vss
c39 78 Vss 3.75522e-19
c40 77 Vss 0.00393043f
c41 72 Vss 0.00270228f
c42 70 Vss 0.00561311f
c43 65 Vss 8.24085e-19
c44 64 Vss 0.0017807f
c45 60 Vss 6.37548e-19
c46 59 Vss 0.00469222f
c47 50 Vss 0.0049931f
c48 41 Vss 7.10513e-22
c49 36 Vss 9.67354e-19
c50 31 Vss 0.00128167f
c51 28 Vss 0.00379689f
c52 23 Vss 0.00389355f
c53 18 Vss 0.089404f
c54 4 Vss 0.134687f
r55 77 80 0.326018
r56 76 77 4.58464
r57 72 76 0.655813
r58 71 78 0.494161
r59 70 80 0.326018
r60 70 71 10.1279
r61 66 78 0.128424
r62 64 78 0.494161
r63 64 65 4.37625
r64 59 65 0.652036
r65 58 60 0.655813
r66 58 59 15.5878
r67 41 72 1.82344
r68 36 50 1.16709
r69 36 66 2.16729
r70 31 60 1.82344
r71 28 41 1.16709
r72 23 31 1.16709
r73 16 50 0.0476429
r74 16 18 2.04225
r75 12 18 0.0685365
r76 6 28 0.185659
r77 4 12 3.8511
r78 2 23 0.185659
.ends

.subckt PM_G2_NOR2_N2_VDD 2 4 6 8 10 27 36 41 45 47 48 52 54 55 58 60 62 64 66
+ 72 78 Vss
c46 78 Vss 0.00511378f
c47 72 Vss 0.00477413f
c48 64 Vss 4.52364e-19
c49 62 Vss 0.00103884f
c50 60 Vss 6.08701e-19
c51 58 Vss 0.00137825f
c52 55 Vss 8.64106e-19
c53 54 Vss 0.00550218f
c54 52 Vss 0.00179763f
c55 49 Vss 0.00174038f
c56 48 Vss 0.00493553f
c57 47 Vss 0.00222713f
c58 45 Vss 0.00953092f
c59 41 Vss 0.00392881f
c60 37 Vss 0.129157f
c61 36 Vss 9.07184e-20
c62 27 Vss 0.035607f
c63 26 Vss 0.102409f
c64 10 Vss 0.13639f
c65 8 Vss 0.134351f
c66 4 Vss 0.13615f
c67 2 Vss 0.137207f
r68 72 75 0.05
r69 62 78 1.16709
r70 60 66 0.326018
r71 60 62 2.16729
r72 58 75 1.16709
r73 56 58 2.20896
r74 54 66 0.326018
r75 54 55 10.1696
r76 50 64 0.0828784
r77 50 52 1.82344
r78 48 56 0.652036
r79 48 49 4.37625
r80 47 55 0.652036
r81 46 64 0.551426
r82 46 47 4.58464
r83 45 64 0.551426
r84 44 49 0.652036
r85 44 45 15.5878
r86 41 52 1.16709
r87 36 72 0.0238214
r88 36 37 2.26917
r89 33 36 2.26917
r90 29 78 0.0476429
r91 27 29 1.5171
r92 26 30 0.652036
r93 26 29 1.4004
r94 23 27 0.652036
r95 20 37 0.00605528
r96 17 33 0.00605528
r97 10 30 3.8511
r98 8 23 3.8511
r99 6 41 0.185659
r100 4 17 3.8511
r101 2 20 3.8511
.ends

.subckt PM_G2_NOR2_N2_B 2 4 10 13 18 21 26 31 Vss
c20 31 Vss 0.00178268f
c21 26 Vss 0.00362926f
c22 18 Vss 0.00103738f
c23 13 Vss 0.112032f
c24 10 Vss 1.01432e-19
c25 2 Vss 0.112208f
r26 23 31 1.16709
r27 21 23 2.04225
r28 18 26 1.16709
r29 18 21 2.79246
r30 13 31 0.50025
r31 10 26 0.50025
r32 4 13 3.09255
r33 2 10 3.09255
.ends

.subckt PM_G2_NOR2_N2_Z 2 4 6 18 22 25 28 Vss
c24 25 Vss 0.00351292f
c25 22 Vss 0.00573209f
c26 18 Vss 0.00386958f
c27 6 Vss 0.00143442f
r28 28 30 4.0845
r29 25 28 6.91864
r30 22 30 1.16709
r31 18 25 1.16709
r32 6 22 0.185659
r33 4 22 0.185659
r34 2 18 0.185659
.ends

.subckt PM_G2_NOR2_N2_A 2 4 10 11 14 18 21 Vss
c17 18 Vss 2.58909e-19
c18 14 Vss 0.170846f
c19 11 Vss 0.0348505f
c20 10 Vss 0.277806f
c21 2 Vss 0.198918f
r22 18 27 1.16709
r23 18 21 0.0416786
r24 14 27 0.05
r25 12 14 1.6338
r26 10 12 0.652036
r27 10 11 8.92755
r28 7 11 0.652036
r29 4 14 4.3179
r30 2 7 5.9517
.ends

.subckt G2_NOR2_N2  VSS VDD B Z A
*
* A	A
* Z	Z
* B	B
* VDD	VDD
* VSS	VSS
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_B_XI3.X0_CG N_VDD_XI3.X0_PGS
+ N_VSS_XI3.X0_S TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VSS_XI4.X0_PGD N_B_XI4.X0_CG N_A_XI4.X0_PGS N_VDD_XI4.X0_S
+ TIGFET_HPNW8
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_VDD_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW8
*
x_PM_G2_NOR2_N2_VSS N_VSS_XI3.X0_S N_VSS_XI4.X0_PGD N_VSS_XI5.X0_S N_VSS_c_2_p
+ N_VSS_c_8_p N_VSS_c_31_p N_VSS_c_3_p N_VSS_c_6_p N_VSS_c_32_p N_VSS_c_13_p
+ N_VSS_c_4_p N_VSS_c_5_p N_VSS_c_14_p N_VSS_c_17_p N_VSS_c_15_p N_VSS_c_20_p
+ N_VSS_c_16_p VSS Vss PM_G2_NOR2_N2_VSS
x_PM_G2_NOR2_N2_VDD N_VDD_XI3.X0_PGD N_VDD_XI3.X0_PGS N_VDD_XI4.X0_S
+ N_VDD_XI5.X0_PGD N_VDD_XI5.X0_PGS N_VDD_c_41_n N_VDD_c_63_p N_VDD_c_71_p
+ N_VDD_c_42_n N_VDD_c_45_n N_VDD_c_47_n N_VDD_c_49_n N_VDD_c_50_n N_VDD_c_56_n
+ N_VDD_c_65_p N_VDD_c_57_n N_VDD_c_58_n N_VDD_c_60_n VDD N_VDD_c_66_p
+ N_VDD_c_61_n Vss PM_G2_NOR2_N2_VDD
x_PM_G2_NOR2_N2_B N_B_XI3.X0_CG N_B_XI4.X0_CG N_B_c_91_n N_B_c_102_p N_B_c_86_n
+ B N_B_c_95_n N_B_c_89_n Vss PM_G2_NOR2_N2_B
x_PM_G2_NOR2_N2_Z N_Z_XI3.X0_D N_Z_XI4.X0_D N_Z_XI5.X0_D N_Z_c_106_n N_Z_c_108_n
+ N_Z_c_110_n Z Vss PM_G2_NOR2_N2_Z
x_PM_G2_NOR2_N2_A N_A_XI4.X0_PGS N_A_XI5.X0_CG N_A_c_130_n N_A_c_133_n
+ N_A_c_135_n N_A_c_137_n A Vss PM_G2_NOR2_N2_A
cc_1 N_VSS_XI4.X0_PGD N_VDD_XI5.X0_PGD 0.00209355f
cc_2 N_VSS_c_2_p N_VDD_c_41_n 0.00209355f
cc_3 N_VSS_c_3_p N_VDD_c_42_n 0.00187494f
cc_4 N_VSS_c_4_p N_VDD_c_42_n 0.00638215f
cc_5 N_VSS_c_5_p N_VDD_c_42_n 0.00189302f
cc_6 N_VSS_c_6_p N_VDD_c_45_n 4.76491e-19
cc_7 N_VSS_c_4_p N_VDD_c_45_n 0.00344537f
cc_8 N_VSS_c_8_p N_VDD_c_47_n 3.4118e-19
cc_9 N_VSS_c_3_p N_VDD_c_47_n 9.64167e-19
cc_10 N_VSS_c_3_p N_VDD_c_49_n 4.54377e-19
cc_11 N_VSS_c_2_p N_VDD_c_50_n 3.66315e-19
cc_12 N_VSS_c_6_p N_VDD_c_50_n 0.00141228f
cc_13 N_VSS_c_13_p N_VDD_c_50_n 0.00114511f
cc_14 N_VSS_c_14_p N_VDD_c_50_n 0.00350144f
cc_15 N_VSS_c_15_p N_VDD_c_50_n 0.00445328f
cc_16 N_VSS_c_16_p N_VDD_c_50_n 7.74609e-19
cc_17 N_VSS_c_17_p N_VDD_c_56_n 0.0010632f
cc_18 N_VSS_c_15_p N_VDD_c_57_n 0.00147105f
cc_19 N_VSS_c_6_p N_VDD_c_58_n 0.00109227f
cc_20 N_VSS_c_20_p N_VDD_c_58_n 3.86251e-19
cc_21 N_VSS_c_4_p N_VDD_c_60_n 0.00116512f
cc_22 N_VSS_c_6_p N_VDD_c_61_n 3.44698e-19
cc_23 N_VSS_c_13_p N_VDD_c_61_n 6.36088e-19
cc_24 N_VSS_c_6_p N_B_c_86_n 5.58916e-19
cc_25 N_VSS_c_13_p N_B_c_86_n 3.52408e-19
cc_26 N_VSS_c_4_p N_B_c_86_n 0.00152314f
cc_27 N_VSS_c_6_p N_B_c_89_n 3.2351e-19
cc_28 N_VSS_c_13_p N_B_c_89_n 0.00119577f
cc_29 N_VSS_c_8_p N_Z_c_106_n 3.43419e-19
cc_30 N_VSS_c_3_p N_Z_c_106_n 3.48267e-19
cc_31 N_VSS_c_31_p N_Z_c_108_n 3.43419e-19
cc_32 N_VSS_c_32_p N_Z_c_108_n 3.48267e-19
cc_33 N_VSS_c_8_p N_Z_c_110_n 3.48267e-19
cc_34 N_VSS_c_31_p N_Z_c_110_n 3.48267e-19
cc_35 N_VSS_c_3_p N_Z_c_110_n 8.54909e-19
cc_36 N_VSS_c_32_p N_Z_c_110_n 5.71987e-19
cc_37 N_VSS_c_4_p N_Z_c_110_n 7.7813e-19
cc_38 N_VSS_c_15_p N_Z_c_110_n 2.40801e-19
cc_39 N_VSS_XI4.X0_PGD N_A_c_130_n 9.55607e-19
cc_40 N_VDD_c_63_p N_B_c_91_n 8.8401e-19
cc_41 N_VDD_c_42_n N_B_c_86_n 0.00264899f
cc_42 N_VDD_c_65_p N_B_c_86_n 5.00177e-19
cc_43 N_VDD_c_66_p N_B_c_86_n 3.55951e-19
cc_44 N_VDD_c_42_n N_B_c_95_n 5.06499e-19
cc_45 N_VDD_c_65_p N_B_c_95_n 3.43988e-19
cc_46 N_VDD_c_66_p N_B_c_95_n 2.75266e-19
cc_47 N_VDD_c_42_n N_B_c_89_n 3.66936e-19
cc_48 N_VDD_c_71_p N_Z_c_108_n 3.43419e-19
cc_49 N_VDD_c_49_n N_Z_c_108_n 3.72199e-19
cc_50 N_VDD_c_50_n N_Z_c_108_n 3.4118e-19
cc_51 N_VDD_c_71_p N_Z_c_110_n 3.48267e-19
cc_52 N_VDD_c_42_n N_Z_c_110_n 9.15147e-19
cc_53 N_VDD_c_49_n N_Z_c_110_n 7.92786e-19
cc_54 N_VDD_c_50_n N_Z_c_110_n 4.80596e-19
cc_55 N_VDD_XI3.X0_PGD N_A_c_130_n 5.1398e-19
cc_56 N_VDD_XI5.X0_PGD N_A_c_130_n 2.51476e-19
cc_57 N_VDD_XI3.X0_PGS N_A_c_133_n 6.75208e-19
cc_58 N_VDD_c_42_n N_A_c_133_n 4.39208e-19
cc_59 N_VDD_c_58_n N_A_c_135_n 3.47446e-19
cc_60 N_VDD_c_61_n N_A_c_135_n 0.00119807f
cc_61 N_VDD_c_58_n N_A_c_137_n 4.24105e-19
cc_62 N_VDD_c_61_n N_A_c_137_n 3.26762e-19
cc_63 N_B_c_86_n N_Z_c_110_n 0.00741085f
cc_64 N_B_c_95_n N_Z_c_110_n 0.0010409f
cc_65 N_B_c_89_n N_Z_c_110_n 9.42705e-19
cc_66 N_B_c_102_p N_A_XI4.X0_PGS 5.00154e-19
cc_67 N_B_c_89_n N_A_XI4.X0_PGS 7.86826e-19
cc_68 N_B_c_95_n N_A_c_130_n 0.00159105f
cc_69 N_B_c_89_n N_A_c_135_n 7.50183e-19
cc_70 N_Z_c_108_n N_A_c_130_n 4.45882e-19
cc_71 N_Z_c_110_n N_A_c_130_n 9.61158e-19
cc_72 N_Z_c_110_n N_A_c_135_n 0.00108982f
cc_73 N_Z_c_110_n N_A_c_137_n 0.00155484f
*
.ends
*
*
.subckt NOR2_HPNW8 A B Y VDD VSS
xgate (VSS VDD B Y A) G2_NOR2_N2
.ends
*
* File: G2_OAI21_N2.pex.netlist
* Created: Wed Mar  2 11:29:59 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_OAI21_N2_VSS 2 4 6 8 10 22 29 37 42 45 50 55 64 73 74 78 84 86 91
+ 94 Vss
c51 92 Vss 5.73928e-19
c52 91 Vss 0.00804514f
c53 86 Vss 0.00176984f
c54 84 Vss 0.00284334f
c55 79 Vss 0.00136792f
c56 78 Vss 0.00717474f
c57 74 Vss 6.26507e-19
c58 73 Vss 0.00636709f
c59 64 Vss 0.0055272f
c60 55 Vss 2.73987e-19
c61 50 Vss 0.00176484f
c62 45 Vss 0.00142483f
c63 42 Vss 0.00389683f
c64 37 Vss 0.00480057f
c65 33 Vss 0.0307649f
c66 29 Vss 6.10339e-20
c67 26 Vss 0.101243f
c68 22 Vss 0.0345703f
c69 21 Vss 0.0712517f
c70 10 Vss 0.136616f
c71 8 Vss 0.135636f
c72 4 Vss 0.135245f
r73 91 94 0.326018
r74 90 91 16.0879
r75 86 90 0.655813
r76 85 92 0.494161
r77 84 94 0.326018
r78 84 85 4.33457
r79 80 92 0.128424
r80 78 92 0.494161
r81 78 79 10.1696
r82 73 79 0.652036
r83 72 74 0.655813
r84 72 73 16.0879
r85 55 86 1.82344
r86 50 64 1.16709
r87 50 80 2.16729
r88 45 74 1.82344
r89 42 55 1.16709
r90 37 45 1.16709
r91 29 64 0.238214
r92 27 33 0.494161
r93 27 29 1.5171
r94 26 30 0.652036
r95 26 29 1.4004
r96 23 33 0.128424
r97 21 33 0.494161
r98 21 22 2.8008
r99 18 22 0.652036
r100 10 30 3.8511
r101 8 23 3.8511
r102 6 42 0.185659
r103 4 18 3.8511
r104 2 37 0.185659
.ends

.subckt PM_G2_OAI21_N2_VDD 2 4 6 8 30 35 38 39 41 43 47 49 51 56 59 65 Vss
c49 65 Vss 0.00587512f
c50 57 Vss 5.34798e-19
c51 56 Vss 0.0102152f
c52 55 Vss 0.00177964f
c53 51 Vss 0.00246273f
c54 49 Vss 0.00378116f
c55 47 Vss 0.00135688f
c56 43 Vss 0.00167028f
c57 41 Vss 8.22855e-19
c58 40 Vss 0.00177964f
c59 39 Vss 0.00981195f
c60 38 Vss 0.0104045f
c61 35 Vss 0.0039168f
c62 30 Vss 0.00399277f
c63 25 Vss 0.0856551f
c64 19 Vss 0.0340946f
c65 18 Vss 0.0688517f
c66 6 Vss 0.137594f
c67 2 Vss 0.137999f
r68 55 59 0.326018
r69 55 56 16.0879
r70 51 56 0.655813
r71 51 53 1.82344
r72 50 57 0.494161
r73 49 59 0.326018
r74 49 50 4.37625
r75 47 65 1.16709
r76 45 57 0.128424
r77 45 47 2.16729
r78 41 43 1.82344
r79 39 57 0.494161
r80 39 40 10.1279
r81 38 41 0.655813
r82 37 40 0.652036
r83 37 38 16.0879
r84 35 53 1.16709
r85 30 43 1.16709
r86 25 65 0.238214
r87 23 25 2.04225
r88 20 23 0.0685365
r89 18 23 0.5835
r90 18 19 2.8008
r91 15 19 0.652036
r92 8 35 0.185659
r93 6 20 3.8511
r94 4 30 0.185659
r95 2 15 3.8511
.ends

.subckt PM_G2_OAI21_N2_B 2 4 13 18 21 26 31 Vss
c21 31 Vss 0.00395418f
c22 26 Vss 0.00337806f
c23 18 Vss 6.82306e-19
c24 13 Vss 0.113634f
c25 10 Vss 1.97908e-19
c26 2 Vss 0.112205f
r27 23 31 1.16709
r28 21 23 1.7505
r29 18 26 1.16709
r30 18 21 3.08421
r31 13 31 0.476429
r32 10 26 0.50025
r33 4 13 3.1509
r34 2 10 3.09255
.ends

.subckt PM_G2_OAI21_N2_A 2 4 13 18 21 26 31 36 44 46 Vss
c41 46 Vss 1.69877e-19
c42 36 Vss 0.00272497f
c43 31 Vss 0.00729791f
c44 26 Vss 0.0034552f
c45 21 Vss 0.00215165f
c46 18 Vss 0.0860045f
c47 13 Vss 5.54498e-20
c48 4 Vss 0.112066f
c49 2 Vss 0.138617f
r50 40 46 0.655813
r51 26 36 1.16709
r52 26 46 4.52212
r53 21 31 1.16709
r54 21 44 0.0416786
r55 21 40 10.8364
r56 18 31 0.238214
r57 15 18 1.92555
r58 13 36 0.50025
r59 7 15 0.0685365
r60 4 13 3.09255
r61 2 7 3.8511
.ends

.subckt PM_G2_OAI21_N2_Z 2 4 6 8 23 27 30 33 Vss
c33 30 Vss 0.0014926f
c34 27 Vss 0.00690919f
c35 23 Vss 0.00596354f
c36 8 Vss 0.00143442f
c37 6 Vss 0.00143442f
r38 33 35 4.20954
r39 30 33 6.79361
r40 27 35 1.16709
r41 23 30 1.16709
r42 8 27 0.185659
r43 6 23 0.185659
r44 4 27 0.185659
r45 2 23 0.185659
.ends

.subckt PM_G2_OAI21_N2_C 2 4 6 13 14 17 24 27 30 Vss
c31 27 Vss 4.25339e-19
c32 24 Vss 0.0812712f
c33 17 Vss 0.202681f
c34 14 Vss 0.0348616f
c35 13 Vss 0.246708f
c36 4 Vss 0.235568f
c37 2 Vss 0.235767f
r38 27 30 0.0833571
r39 23 24 2.04225
r40 20 24 0.0685365
r41 17 27 1.16709
r42 15 23 0.0685365
r43 15 17 2.8008
r44 13 23 0.5835
r45 13 14 8.92755
r46 10 14 0.652036
r47 6 17 4.3179
r48 4 20 7.1187
r49 2 10 7.1187
.ends

.subckt G2_OAI21_N2  VSS VDD B A Z C
*
* C	C
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_B_XI3.X0_CG N_C_XI3.X0_PGS N_VSS_XI3.X0_S
+ TIGFET_HPNW8
XI0.X0 N_Z_XI0.X0_D N_VSS_XI0.X0_PGD N_B_XI0.X0_CG N_A_XI0.X0_PGS N_VDD_XI0.X0_S
+ TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VDD_XI4.X0_PGD N_A_XI4.X0_CG N_C_XI4.X0_PGS N_VSS_XI4.X0_S
+ TIGFET_HPNW8
XI2.X0 N_Z_XI2.X0_D N_VSS_XI2.X0_PGD N_C_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW8
*
x_PM_G2_OAI21_N2_VSS N_VSS_XI3.X0_S N_VSS_XI0.X0_PGD N_VSS_XI4.X0_S
+ N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS N_VSS_c_29_p N_VSS_c_46_p N_VSS_c_1_p
+ N_VSS_c_9_p N_VSS_c_2_p N_VSS_c_21_p N_VSS_c_10_p N_VSS_c_22_p N_VSS_c_3_p
+ N_VSS_c_4_p N_VSS_c_8_p N_VSS_c_12_p N_VSS_c_11_p N_VSS_c_14_p VSS Vss
+ PM_G2_OAI21_N2_VSS
x_PM_G2_OAI21_N2_VDD N_VDD_XI3.X0_PGD N_VDD_XI0.X0_S N_VDD_XI4.X0_PGD
+ N_VDD_XI2.X0_S N_VDD_c_84_p N_VDD_c_85_p N_VDD_c_52_n N_VDD_c_56_n
+ N_VDD_c_57_n N_VDD_c_58_n N_VDD_c_77_p N_VDD_c_60_n N_VDD_c_63_n N_VDD_c_66_n
+ VDD N_VDD_c_74_p Vss PM_G2_OAI21_N2_VDD
x_PM_G2_OAI21_N2_B N_B_XI3.X0_CG N_B_XI0.X0_CG N_B_c_109_p N_B_c_101_n B
+ N_B_c_104_n N_B_c_105_n Vss PM_G2_OAI21_N2_B
x_PM_G2_OAI21_N2_A N_A_XI0.X0_PGS N_A_XI4.X0_CG N_A_c_137_n N_A_c_145_n
+ N_A_c_123_n N_A_c_128_n N_A_c_130_n N_A_c_134_n A N_A_c_135_n Vss
+ PM_G2_OAI21_N2_A
x_PM_G2_OAI21_N2_Z N_Z_XI3.X0_D N_Z_XI0.X0_D N_Z_XI4.X0_D N_Z_XI2.X0_D
+ N_Z_c_163_n N_Z_c_174_n N_Z_c_167_n Z Vss PM_G2_OAI21_N2_Z
x_PM_G2_OAI21_N2_C N_C_XI3.X0_PGS N_C_XI4.X0_PGS N_C_XI2.X0_CG N_C_c_196_n
+ N_C_c_218_n N_C_c_198_n N_C_c_201_n N_C_c_202_n C Vss PM_G2_OAI21_N2_C
cc_1 N_VSS_c_1_p N_VDD_c_52_n 9.5668e-19
cc_2 N_VSS_c_2_p N_VDD_c_52_n 0.00165395f
cc_3 N_VSS_c_3_p N_VDD_c_52_n 0.00691557f
cc_4 N_VSS_c_4_p N_VDD_c_52_n 0.00189413f
cc_5 N_VSS_c_2_p N_VDD_c_56_n 9.07068e-19
cc_6 N_VSS_c_3_p N_VDD_c_57_n 0.0016897f
cc_7 N_VSS_c_2_p N_VDD_c_58_n 4.55601e-19
cc_8 N_VSS_c_8_p N_VDD_c_58_n 4.44911e-19
cc_9 N_VSS_c_9_p N_VDD_c_60_n 3.02646e-19
cc_10 N_VSS_c_10_p N_VDD_c_60_n 4.09912e-19
cc_11 N_VSS_c_11_p N_VDD_c_60_n 4.66923e-19
cc_12 N_VSS_c_12_p N_VDD_c_63_n 4.44911e-19
cc_13 N_VSS_c_11_p N_VDD_c_63_n 4.55601e-19
cc_14 N_VSS_c_14_p N_VDD_c_63_n 0.00176782f
cc_15 N_VSS_c_9_p N_VDD_c_66_n 9.5668e-19
cc_16 N_VSS_c_10_p N_VDD_c_66_n 0.00165395f
cc_17 N_VSS_c_11_p N_VDD_c_66_n 0.00189413f
cc_18 N_VSS_c_14_p N_VDD_c_66_n 0.00744813f
cc_19 N_VSS_c_3_p N_B_c_101_n 5.69535e-19
cc_20 N_VSS_XI0.X0_PGD N_A_XI0.X0_PGS 0.00176902f
cc_21 N_VSS_c_21_p N_A_c_123_n 8.59446e-19
cc_22 N_VSS_c_22_p N_A_c_123_n 3.44698e-19
cc_23 N_VSS_c_3_p N_A_c_123_n 0.003788f
cc_24 N_VSS_c_8_p N_A_c_123_n 0.00211252f
cc_25 N_VSS_c_14_p N_A_c_123_n 0.00180094f
cc_26 N_VSS_c_8_p N_A_c_128_n 7.40806e-19
cc_27 N_VSS_c_14_p N_A_c_128_n 7.9739e-19
cc_28 N_VSS_XI0.X0_PGD N_A_c_130_n 3.11814e-19
cc_29 N_VSS_c_29_p N_A_c_130_n 0.00322564f
cc_30 N_VSS_c_21_p N_A_c_130_n 3.44698e-19
cc_31 N_VSS_c_22_p N_A_c_130_n 6.61253e-19
cc_32 N_VSS_c_22_p N_A_c_134_n 2.86526e-19
cc_33 N_VSS_c_3_p N_A_c_135_n 0.00310102f
cc_34 N_VSS_c_1_p N_Z_c_163_n 3.43419e-19
cc_35 N_VSS_c_9_p N_Z_c_163_n 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_c_163_n 3.48267e-19
cc_37 N_VSS_c_10_p N_Z_c_163_n 3.48267e-19
cc_38 N_VSS_c_1_p N_Z_c_167_n 3.48267e-19
cc_39 N_VSS_c_9_p N_Z_c_167_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_167_n 5.71987e-19
cc_41 N_VSS_c_10_p N_Z_c_167_n 5.71987e-19
cc_42 N_VSS_c_8_p N_Z_c_167_n 3.27942e-19
cc_43 N_VSS_c_14_p N_Z_c_167_n 6.37542e-19
cc_44 N_VSS_XI0.X0_PGD N_C_c_196_n 6.82193e-19
cc_45 N_VSS_XI2.X0_PGD N_C_c_196_n 6.82193e-19
cc_46 N_VSS_c_46_p N_C_c_198_n 4.58946e-19
cc_47 N_VSS_c_21_p N_C_c_198_n 2.87758e-19
cc_48 N_VSS_c_22_p N_C_c_198_n 0.00236077f
cc_49 N_VSS_XI2.X0_PGS N_C_c_201_n 8.15793e-19
cc_50 N_VSS_c_21_p N_C_c_202_n 2.83343e-19
cc_51 N_VSS_c_22_p N_C_c_202_n 2.87758e-19
cc_52 N_VDD_c_52_n N_B_c_101_n 0.00231792f
cc_53 N_VDD_c_56_n N_B_c_101_n 2.08521e-19
cc_54 N_VDD_c_52_n N_B_c_104_n 3.66936e-19
cc_55 N_VDD_c_52_n N_B_c_105_n 4.5927e-19
cc_56 N_VDD_c_74_p N_A_XI4.X0_CG 0.00253477f
cc_57 N_VDD_c_74_p N_A_c_137_n 6.39343e-19
cc_58 N_VDD_c_56_n N_A_c_128_n 7.76297e-19
cc_59 N_VDD_c_77_p N_A_c_128_n 5.10019e-19
cc_60 N_VDD_c_66_n N_A_c_128_n 6.23587e-19
cc_61 N_VDD_c_74_p N_A_c_128_n 3.18657e-19
cc_62 N_VDD_c_66_n N_A_c_134_n 3.66936e-19
cc_63 N_VDD_c_74_p N_A_c_134_n 6.82215e-19
cc_64 N_VDD_c_52_n N_A_c_135_n 6.11072e-19
cc_65 N_VDD_c_56_n N_Z_c_163_n 3.02646e-19
cc_66 N_VDD_c_84_p N_Z_c_174_n 3.43419e-19
cc_67 N_VDD_c_85_p N_Z_c_174_n 3.43419e-19
cc_68 N_VDD_c_58_n N_Z_c_174_n 3.72199e-19
cc_69 N_VDD_c_63_n N_Z_c_174_n 3.72199e-19
cc_70 N_VDD_c_84_p N_Z_c_167_n 3.48267e-19
cc_71 N_VDD_c_85_p N_Z_c_167_n 3.48267e-19
cc_72 N_VDD_c_52_n N_Z_c_167_n 7.99049e-19
cc_73 N_VDD_c_56_n N_Z_c_167_n 6.12187e-19
cc_74 N_VDD_c_58_n N_Z_c_167_n 5.09542e-19
cc_75 N_VDD_c_63_n N_Z_c_167_n 7.72285e-19
cc_76 N_VDD_c_66_n N_Z_c_167_n 0.00141871f
cc_77 N_VDD_c_52_n N_C_XI3.X0_PGS 6.13097e-19
cc_78 N_VDD_c_66_n N_C_XI4.X0_PGS 6.32546e-19
cc_79 N_VDD_XI3.X0_PGD N_C_c_196_n 6.82193e-19
cc_80 N_VDD_XI4.X0_PGD N_C_c_196_n 6.82193e-19
cc_81 N_VDD_c_66_n N_C_c_198_n 5.55044e-19
cc_82 N_VDD_c_66_n N_C_c_202_n 5.04211e-19
cc_83 N_B_c_105_n N_A_c_145_n 4.64013e-19
cc_84 N_B_c_101_n N_A_c_123_n 0.0028587f
cc_85 N_B_c_105_n N_A_c_123_n 2.87758e-19
cc_86 N_B_c_109_p N_A_c_130_n 0.00249847f
cc_87 N_B_c_101_n N_A_c_130_n 3.4348e-19
cc_88 N_B_c_105_n N_A_c_130_n 6.82215e-19
cc_89 N_B_c_104_n N_A_c_134_n 8.86454e-19
cc_90 N_B_c_101_n N_A_c_135_n 7.33011e-19
cc_91 N_B_c_101_n N_Z_c_167_n 0.00671f
cc_92 N_B_c_104_n N_Z_c_167_n 9.58174e-19
cc_93 N_B_c_105_n N_Z_c_167_n 0.00100281f
cc_94 N_B_XI3.X0_CG N_C_XI3.X0_PGS 4.87172e-19
cc_95 N_B_c_104_n N_C_XI3.X0_PGS 0.001089f
cc_96 N_B_c_104_n N_C_c_196_n 6.02551e-19
cc_97 N_B_c_105_n N_C_c_196_n 0.00129343f
cc_98 N_B_c_105_n N_C_c_198_n 9.54365e-19
cc_99 N_A_c_123_n N_Z_c_167_n 0.00174866f
cc_100 N_A_c_128_n N_Z_c_167_n 0.00351012f
cc_101 N_A_c_134_n N_Z_c_167_n 9.53427e-19
cc_102 N_A_XI4.X0_CG N_C_XI4.X0_PGS 4.87172e-19
cc_103 N_A_c_134_n N_C_XI4.X0_PGS 0.001089f
cc_104 N_A_c_134_n N_C_c_196_n 0.00151445f
cc_105 N_A_XI0.X0_PGS N_C_c_218_n 8.15793e-19
cc_106 N_A_c_128_n N_C_c_198_n 5.38228e-19
cc_107 N_A_c_134_n N_C_c_198_n 0.00209031f
cc_108 N_A_c_128_n N_C_c_202_n 8.16123e-19
cc_109 N_Z_c_163_n N_C_c_196_n 3.50149e-19
cc_110 N_Z_c_174_n N_C_c_196_n 3.50149e-19
cc_111 N_Z_c_167_n N_C_c_196_n 3.56555e-19
cc_112 N_Z_c_167_n N_C_c_198_n 0.00102535f
cc_113 N_Z_c_167_n N_C_c_202_n 0.00141616f
*
.ends
*
*
.subckt OAI21_HPNW8 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 A0 Y B0) G2_OAI21_N2
.ends
*
* File: G3_OR2_N2.pex.netlist
* Created: Tue Mar  1 12:00:05 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_OR2_N2_VSS 2 4 6 8 10 12 28 29 38 44 49 52 57 62 67 76 85 90 91 93
+ 97 98 103 109 115 116 Vss
c69 116 Vss 3.88979e-19
c70 115 Vss 3.75522e-19
c71 109 Vss 0.00356171f
c72 103 Vss 0.00288176f
c73 98 Vss 8.31407e-19
c74 97 Vss 0.0017807f
c75 91 Vss 6.38539e-19
c76 90 Vss 0.00489715f
c77 85 Vss 0.00399322f
c78 76 Vss 0.00493786f
c79 67 Vss 5.89061e-19
c80 62 Vss 7.90818e-19
c81 57 Vss 8.66334e-19
c82 52 Vss 0.00128155f
c83 49 Vss 0.00709351f
c84 44 Vss 0.00389355f
c85 38 Vss 0.0895618f
c86 29 Vss 0.0349332f
c87 28 Vss 0.0997249f
c88 12 Vss 0.134814f
c89 10 Vss 0.13405f
c90 8 Vss 0.00143442f
c91 4 Vss 0.134687f
r92 110 116 0.494161
r93 109 111 0.652036
r94 109 110 7.46046
r95 105 116 0.128424
r96 104 115 0.494161
r97 103 116 0.494161
r98 103 104 7.46046
r99 99 115 0.128424
r100 97 115 0.494161
r101 97 98 4.37625
r102 91 93 0.765844
r103 90 98 0.652036
r104 89 91 0.655813
r105 89 90 15.5878
r106 67 85 1.16709
r107 67 111 2.16729
r108 62 105 5.2515
r109 57 76 1.16709
r110 57 99 2.16729
r111 52 93 1.05759
r112 49 62 1.16709
r113 44 52 1.16709
r114 36 76 0.0476429
r115 36 38 2.04225
r116 31 85 0.0476429
r117 29 31 1.45875
r118 28 32 0.652036
r119 28 31 1.45875
r120 25 29 0.652036
r121 22 38 0.0685365
r122 12 32 3.8511
r123 10 25 3.8511
r124 8 49 0.185659
r125 6 49 0.185659
r126 4 22 3.8511
r127 2 44 0.185659
.ends

.subckt PM_G3_OR2_N2_VDD 2 4 6 8 10 12 14 16 37 46 56 62 67 70 72 73 77 79 80 83
+ 87 89 93 95 97 102 104 105 106 107 113 119 124 Vss
c78 124 Vss 0.00436477f
c79 119 Vss 0.00478009f
c80 113 Vss 0.00477414f
c81 107 Vss 2.39889e-19
c82 106 Vss 2.39889e-19
c83 105 Vss 4.52364e-19
c84 102 Vss 0.00334204f
c85 97 Vss 0.00329381f
c86 95 Vss 0.00842218f
c87 93 Vss 5.48147e-19
c88 89 Vss 0.00206676f
c89 87 Vss 4.88586e-19
c90 83 Vss 0.00135406f
c91 80 Vss 8.68155e-19
c92 79 Vss 0.00563376f
c93 77 Vss 0.0017975f
c94 73 Vss 0.0049339f
c95 72 Vss 0.00221679f
c96 70 Vss 0.00947695f
c97 69 Vss 0.00174028f
c98 67 Vss 0.00532741f
c99 62 Vss 0.00393183f
c100 57 Vss 0.129157f
c101 56 Vss 9.10906e-20
c102 47 Vss 0.0358563f
c103 46 Vss 0.101295f
c104 37 Vss 0.035607f
c105 36 Vss 0.101546f
c106 14 Vss 0.134527f
c107 12 Vss 0.134502f
c108 10 Vss 0.13477f
c109 8 Vss 0.134351f
c110 4 Vss 0.136655f
c111 2 Vss 0.137748f
r112 113 116 0.05
r113 101 102 4.58464
r114 97 101 0.655813
r115 97 99 1.82344
r116 96 107 0.494161
r117 95 102 0.652036
r118 95 96 10.1279
r119 93 124 1.16709
r120 91 107 0.128424
r121 91 93 2.16729
r122 90 106 0.494161
r123 89 107 0.494161
r124 89 90 4.54296
r125 87 119 1.16709
r126 85 106 0.128424
r127 85 87 2.16729
r128 83 116 1.16709
r129 81 83 2.16729
r130 79 106 0.494161
r131 79 80 10.1696
r132 75 105 0.0828784
r133 75 77 1.82344
r134 74 104 0.326018
r135 73 81 0.652036
r136 73 74 4.37625
r137 72 80 0.652036
r138 71 105 0.551426
r139 71 72 4.58464
r140 70 105 0.551426
r141 69 104 0.326018
r142 69 70 15.5461
r143 67 99 1.16709
r144 62 77 1.16709
r145 56 113 0.0238214
r146 56 57 2.26917
r147 53 56 2.26917
r148 49 124 0.0476429
r149 47 49 1.45875
r150 46 50 0.652036
r151 46 49 1.45875
r152 43 47 0.652036
r153 39 119 0.0476429
r154 37 39 1.5171
r155 36 40 0.652036
r156 36 39 1.4004
r157 33 37 0.652036
r158 30 57 0.00605528
r159 27 53 0.00605528
r160 16 67 0.185659
r161 14 43 3.8511
r162 12 50 3.8511
r163 10 40 3.8511
r164 8 33 3.8511
r165 6 62 0.185659
r166 4 27 3.8511
r167 2 30 3.8511
.ends

.subckt PM_G3_OR2_N2_B 2 4 10 13 18 21 26 31 Vss
c21 31 Vss 0.00178268f
c22 26 Vss 0.00362926f
c23 18 Vss 9.47382e-19
c24 13 Vss 0.112032f
c25 10 Vss 1.01848e-19
c26 2 Vss 0.112208f
r27 23 31 1.16709
r28 21 23 2.20896
r29 18 26 1.16709
r30 18 21 2.62575
r31 13 31 0.50025
r32 10 26 0.50025
r33 4 13 3.09255
r34 2 10 3.09255
.ends

.subckt PM_G3_OR2_N2_NET21 2 4 6 8 10 24 27 38 42 45 53 66 70 Vss
c39 70 Vss 0.00743392f
c40 66 Vss 0.0057739f
c41 53 Vss 0.00155523f
c42 45 Vss 0.00308587f
c43 42 Vss 0.00569159f
c44 38 Vss 0.00386958f
c45 27 Vss 1.05421e-19
c46 24 Vss 0.225855f
c47 21 Vss 0.125908f
c48 19 Vss 0.0247918f
c49 10 Vss 0.139046f
c50 6 Vss 0.00143442f
r51 70 74 0.655813
r52 53 66 1.16709
r53 53 74 2.08393
r54 48 70 7.03847
r55 48 50 5.835
r56 45 48 5.16814
r57 42 50 1.16709
r58 38 45 1.16709
r59 27 66 0.0476429
r60 25 27 0.326018
r61 25 27 0.1167
r62 24 28 0.652036
r63 24 27 6.7686
r64 21 66 0.357321
r65 19 27 0.326018
r66 19 21 0.40845
r67 10 28 3.8511
r68 8 21 3.44265
r69 6 42 0.185659
r70 4 42 0.185659
r71 2 38 0.185659
.ends

.subckt PM_G3_OR2_N2_A 2 4 10 11 14 18 21 Vss
c21 18 Vss 3.18373e-19
c22 14 Vss 0.170625f
c23 11 Vss 0.0348505f
c24 10 Vss 0.277805f
c25 2 Vss 0.198918f
r26 18 27 1.16709
r27 18 21 0.0833571
r28 14 27 0.05
r29 12 14 1.6338
r30 10 12 0.652036
r31 10 11 8.92755
r32 7 11 0.652036
r33 4 14 4.3179
r34 2 7 5.9517
.ends

.subckt PM_G3_OR2_N2_Z 2 4 13 16 19 Vss
c12 13 Vss 0.00522942f
c13 4 Vss 0.00143442f
r14 16 19 0.0353636
r15 13 19 1.16709
r16 4 13 0.185659
r17 2 13 0.185659
.ends

.subckt G3_OR2_N2  VSS VDD B A Z
*
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI7.X0 N_NET21_XI7.X0_D N_VDD_XI7.X0_PGD N_B_XI7.X0_CG N_VDD_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW8
XI5.X0 N_NET21_XI5.X0_D N_VSS_XI5.X0_PGD N_B_XI5.X0_CG N_A_XI5.X0_PGS
+ N_VDD_XI5.X0_S TIGFET_HPNW8
XI6.X0 N_NET21_XI6.X0_D N_VDD_XI6.X0_PGD N_A_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW8
XI8.X0 N_Z_XI8.X0_D N_VDD_XI8.X0_PGD N_NET21_XI8.X0_CG N_VDD_XI8.X0_PGS
+ N_VSS_XI8.X0_S TIGFET_HPNW8
XI9.X0 N_Z_XI9.X0_D N_VSS_XI9.X0_PGD N_NET21_XI9.X0_CG N_VSS_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW8
*
x_PM_G3_OR2_N2_VSS N_VSS_XI7.X0_S N_VSS_XI5.X0_PGD N_VSS_XI6.X0_S N_VSS_XI8.X0_S
+ N_VSS_XI9.X0_PGD N_VSS_XI9.X0_PGS N_VSS_c_30_p N_VSS_c_4_p N_VSS_c_3_p
+ N_VSS_c_10_p N_VSS_c_53_p N_VSS_c_5_p N_VSS_c_8_p N_VSS_c_21_p N_VSS_c_28_p
+ N_VSS_c_15_p N_VSS_c_29_p N_VSS_c_6_p N_VSS_c_7_p VSS N_VSS_c_16_p
+ N_VSS_c_19_p N_VSS_c_17_p N_VSS_c_25_p N_VSS_c_18_p N_VSS_c_26_p Vss
+ PM_G3_OR2_N2_VSS
x_PM_G3_OR2_N2_VDD N_VDD_XI7.X0_PGD N_VDD_XI7.X0_PGS N_VDD_XI5.X0_S
+ N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI8.X0_PGD N_VDD_XI8.X0_PGS
+ N_VDD_XI9.X0_S N_VDD_c_72_n N_VDD_c_73_n N_VDD_c_114_p N_VDD_c_124_p
+ N_VDD_c_142_p N_VDD_c_74_n N_VDD_c_77_n N_VDD_c_79_n N_VDD_c_81_n N_VDD_c_82_n
+ N_VDD_c_88_n N_VDD_c_116_p N_VDD_c_89_n N_VDD_c_92_n N_VDD_c_96_n N_VDD_c_99_n
+ N_VDD_c_144_p N_VDD_c_104_n VDD N_VDD_c_107_n N_VDD_c_108_n N_VDD_c_109_n
+ N_VDD_c_117_p N_VDD_c_110_n N_VDD_c_112_n Vss PM_G3_OR2_N2_VDD
x_PM_G3_OR2_N2_B N_B_XI7.X0_CG N_B_XI5.X0_CG N_B_c_153_n N_B_c_165_p N_B_c_148_n
+ B N_B_c_157_n N_B_c_151_n Vss PM_G3_OR2_N2_B
x_PM_G3_OR2_N2_NET21 N_NET21_XI7.X0_D N_NET21_XI5.X0_D N_NET21_XI6.X0_D
+ N_NET21_XI8.X0_CG N_NET21_XI9.X0_CG N_NET21_c_169_n N_NET21_c_184_n
+ N_NET21_c_170_n N_NET21_c_172_n N_NET21_c_174_n N_NET21_c_179_n
+ N_NET21_c_194_n N_NET21_c_180_n Vss PM_G3_OR2_N2_NET21
x_PM_G3_OR2_N2_A N_A_XI5.X0_PGS N_A_XI6.X0_CG N_A_c_208_n N_A_c_211_n
+ N_A_c_213_n N_A_c_215_n A Vss PM_G3_OR2_N2_A
x_PM_G3_OR2_N2_Z N_Z_XI8.X0_D N_Z_XI9.X0_D N_Z_c_229_n Z N_Z_c_231_n Vss
+ PM_G3_OR2_N2_Z
cc_1 N_VSS_XI5.X0_PGD N_VDD_XI6.X0_PGD 0.00204282f
cc_2 N_VSS_XI9.X0_PGD N_VDD_XI8.X0_PGD 0.00196484f
cc_3 N_VSS_c_3_p N_VDD_c_72_n 0.00204282f
cc_4 N_VSS_c_4_p N_VDD_c_73_n 0.00196484f
cc_5 N_VSS_c_5_p N_VDD_c_74_n 0.00187494f
cc_6 N_VSS_c_6_p N_VDD_c_74_n 0.00677253f
cc_7 N_VSS_c_7_p N_VDD_c_74_n 0.00189302f
cc_8 N_VSS_c_8_p N_VDD_c_77_n 4.76491e-19
cc_9 N_VSS_c_6_p N_VDD_c_77_n 0.0033599f
cc_10 N_VSS_c_10_p N_VDD_c_79_n 3.44698e-19
cc_11 N_VSS_c_5_p N_VDD_c_79_n 9.72065e-19
cc_12 N_VSS_c_5_p N_VDD_c_81_n 4.54347e-19
cc_13 N_VSS_c_3_p N_VDD_c_82_n 3.66315e-19
cc_14 N_VSS_c_8_p N_VDD_c_82_n 0.00141228f
cc_15 N_VSS_c_15_p N_VDD_c_82_n 0.00114511f
cc_16 N_VSS_c_16_p N_VDD_c_82_n 0.00350144f
cc_17 N_VSS_c_17_p N_VDD_c_82_n 0.00435073f
cc_18 N_VSS_c_18_p N_VDD_c_82_n 7.74609e-19
cc_19 N_VSS_c_19_p N_VDD_c_88_n 0.00106851f
cc_20 N_VSS_c_8_p N_VDD_c_89_n 8.39054e-19
cc_21 N_VSS_c_21_p N_VDD_c_89_n 3.93845e-19
cc_22 N_VSS_c_15_p N_VDD_c_89_n 3.95933e-19
cc_23 N_VSS_c_21_p N_VDD_c_92_n 4.34701e-19
cc_24 N_VSS_c_17_p N_VDD_c_92_n 0.00137965f
cc_25 N_VSS_c_25_p N_VDD_c_92_n 0.00142692f
cc_26 N_VSS_c_26_p N_VDD_c_92_n 0.00107375f
cc_27 N_VSS_c_21_p N_VDD_c_96_n 3.91951e-19
cc_28 N_VSS_c_28_p N_VDD_c_96_n 8.45954e-19
cc_29 N_VSS_c_29_p N_VDD_c_96_n 3.99794e-19
cc_30 N_VSS_c_30_p N_VDD_c_99_n 4.1253e-19
cc_31 N_VSS_c_4_p N_VDD_c_99_n 3.9313e-19
cc_32 N_VSS_c_28_p N_VDD_c_99_n 0.00161703f
cc_33 N_VSS_c_29_p N_VDD_c_99_n 2.26455e-19
cc_34 N_VSS_c_25_p N_VDD_c_99_n 0.00609002f
cc_35 N_VSS_XI9.X0_PGS N_VDD_c_104_n 3.05236e-19
cc_36 N_VSS_c_28_p N_VDD_c_104_n 8.67538e-19
cc_37 N_VSS_c_29_p N_VDD_c_104_n 3.66936e-19
cc_38 N_VSS_c_6_p N_VDD_c_107_n 0.00116512f
cc_39 N_VSS_c_17_p N_VDD_c_108_n 9.95024e-19
cc_40 N_VSS_c_25_p N_VDD_c_109_n 9.97484e-19
cc_41 N_VSS_c_8_p N_VDD_c_110_n 3.44698e-19
cc_42 N_VSS_c_15_p N_VDD_c_110_n 6.36088e-19
cc_43 N_VSS_c_28_p N_VDD_c_112_n 3.48267e-19
cc_44 N_VSS_c_29_p N_VDD_c_112_n 6.489e-19
cc_45 N_VSS_c_8_p N_B_c_148_n 5.58916e-19
cc_46 N_VSS_c_15_p N_B_c_148_n 3.52408e-19
cc_47 N_VSS_c_6_p N_B_c_148_n 8.9847e-19
cc_48 N_VSS_c_8_p N_B_c_151_n 3.2351e-19
cc_49 N_VSS_c_15_p N_B_c_151_n 0.00119577f
cc_50 N_VSS_XI9.X0_PGD N_NET21_c_169_n 4.25712e-19
cc_51 N_VSS_c_10_p N_NET21_c_170_n 3.43419e-19
cc_52 N_VSS_c_5_p N_NET21_c_170_n 3.48267e-19
cc_53 N_VSS_c_53_p N_NET21_c_172_n 3.43419e-19
cc_54 N_VSS_c_21_p N_NET21_c_172_n 3.48267e-19
cc_55 N_VSS_c_10_p N_NET21_c_174_n 3.48267e-19
cc_56 N_VSS_c_53_p N_NET21_c_174_n 3.48267e-19
cc_57 N_VSS_c_5_p N_NET21_c_174_n 8.54909e-19
cc_58 N_VSS_c_21_p N_NET21_c_174_n 5.71987e-19
cc_59 N_VSS_c_6_p N_NET21_c_174_n 6.84771e-19
cc_60 N_VSS_c_25_p N_NET21_c_179_n 2.36784e-19
cc_61 N_VSS_c_21_p N_NET21_c_180_n 9.51297e-19
cc_62 N_VSS_c_6_p N_NET21_c_180_n 2.32409e-19
cc_63 N_VSS_c_17_p N_NET21_c_180_n 8.71002e-19
cc_64 N_VSS_XI5.X0_PGD N_A_c_208_n 9.55607e-19
cc_65 N_VSS_c_53_p N_Z_c_229_n 3.43419e-19
cc_66 N_VSS_c_21_p N_Z_c_229_n 3.48267e-19
cc_67 N_VSS_c_53_p N_Z_c_231_n 3.48267e-19
cc_68 N_VSS_c_21_p N_Z_c_231_n 7.85754e-19
cc_69 N_VSS_c_25_p N_Z_c_231_n 2.50289e-19
cc_70 N_VDD_c_114_p N_B_c_153_n 8.95172e-19
cc_71 N_VDD_c_74_n N_B_c_148_n 0.00268777f
cc_72 N_VDD_c_116_p N_B_c_148_n 5.04982e-19
cc_73 N_VDD_c_117_p N_B_c_148_n 3.55951e-19
cc_74 N_VDD_c_74_n N_B_c_157_n 5.06499e-19
cc_75 N_VDD_c_116_p N_B_c_157_n 3.47446e-19
cc_76 N_VDD_c_117_p N_B_c_157_n 2.75266e-19
cc_77 N_VDD_c_74_n N_B_c_151_n 3.66936e-19
cc_78 N_VDD_XI8.X0_PGD N_NET21_c_169_n 4.28909e-19
cc_79 N_VDD_c_112_n N_NET21_c_184_n 9.53212e-19
cc_80 N_VDD_c_124_p N_NET21_c_172_n 3.43419e-19
cc_81 N_VDD_c_81_n N_NET21_c_172_n 3.72199e-19
cc_82 N_VDD_c_82_n N_NET21_c_172_n 3.4118e-19
cc_83 N_VDD_c_124_p N_NET21_c_174_n 3.48267e-19
cc_84 N_VDD_c_74_n N_NET21_c_174_n 8.27149e-19
cc_85 N_VDD_c_81_n N_NET21_c_174_n 7.92786e-19
cc_86 N_VDD_c_82_n N_NET21_c_174_n 4.80596e-19
cc_87 N_VDD_c_96_n N_NET21_c_179_n 3.42685e-19
cc_88 N_VDD_c_112_n N_NET21_c_179_n 3.2351e-19
cc_89 N_VDD_c_112_n N_NET21_c_194_n 2.68747e-19
cc_90 N_VDD_XI7.X0_PGD N_A_c_208_n 5.1398e-19
cc_91 N_VDD_XI6.X0_PGD N_A_c_208_n 2.51476e-19
cc_92 N_VDD_XI7.X0_PGS N_A_c_211_n 6.75208e-19
cc_93 N_VDD_c_74_n N_A_c_211_n 4.39208e-19
cc_94 N_VDD_c_89_n N_A_c_213_n 3.47446e-19
cc_95 N_VDD_c_110_n N_A_c_213_n 0.00119807f
cc_96 N_VDD_c_89_n N_A_c_215_n 4.0116e-19
cc_97 N_VDD_c_110_n N_A_c_215_n 3.26762e-19
cc_98 N_VDD_c_142_p N_Z_c_229_n 3.43419e-19
cc_99 N_VDD_c_99_n N_Z_c_229_n 3.4118e-19
cc_100 N_VDD_c_144_p N_Z_c_229_n 3.72199e-19
cc_101 N_VDD_c_142_p N_Z_c_231_n 3.48267e-19
cc_102 N_VDD_c_99_n N_Z_c_231_n 4.63968e-19
cc_103 N_VDD_c_144_p N_Z_c_231_n 7.4527e-19
cc_104 N_B_c_148_n N_NET21_c_174_n 0.00749505f
cc_105 N_B_c_157_n N_NET21_c_174_n 0.0010409f
cc_106 N_B_c_151_n N_NET21_c_174_n 9.42705e-19
cc_107 N_B_c_148_n N_NET21_c_180_n 2.06853e-19
cc_108 N_B_c_165_p N_A_XI5.X0_PGS 5.00154e-19
cc_109 N_B_c_151_n N_A_XI5.X0_PGS 7.86826e-19
cc_110 N_B_c_157_n N_A_c_208_n 0.0015904f
cc_111 N_B_c_151_n N_A_c_213_n 7.50183e-19
cc_112 N_NET21_c_172_n N_A_c_208_n 4.45882e-19
cc_113 N_NET21_c_174_n N_A_c_208_n 8.51551e-19
cc_114 N_NET21_c_174_n N_A_c_213_n 0.00108501f
cc_115 N_NET21_c_179_n N_A_c_213_n 3.48267e-19
cc_116 N_NET21_c_194_n N_A_c_213_n 0.00171208f
cc_117 N_NET21_c_174_n N_A_c_215_n 0.0014331f
cc_118 N_NET21_c_179_n N_A_c_215_n 4.16154e-19
cc_119 N_NET21_c_180_n N_A_c_215_n 3.53251e-19
cc_120 N_NET21_c_169_n N_Z_c_229_n 6.55689e-19
*
.ends
*
*
.subckt OR2_HPNW8 A B Y VDD VSS
xgate (VSS VDD B A Y) G3_OR2_N2
.ends
*
* File: G4_XNOR2_N2.pex.netlist
* Created: Wed Mar 16 11:10:33 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XNOR2_N2_VDD 2 5 9 12 14 16 32 42 43 45 54 59 63 66 68 69 70 73 75
+ 76 79 81 85 89 91 93 98 99 100 103 109 114 Vss
c104 114 Vss 0.00451172f
c105 109 Vss 0.0046333f
c106 101 Vss 8.60971e-19
c107 100 Vss 2.39889e-19
c108 99 Vss 4.52364e-19
c109 98 Vss 0.00501239f
c110 93 Vss 0.00287584f
c111 91 Vss 0.0106993f
c112 89 Vss 0.00158164f
c113 85 Vss 4.92677e-19
c114 81 Vss 0.00450584f
c115 79 Vss 0.00110794f
c116 76 Vss 8.67986e-19
c117 75 Vss 0.00221168f
c118 73 Vss 0.00195091f
c119 70 Vss 8.63914e-19
c120 69 Vss 0.005504f
c121 68 Vss 0.00838153f
c122 66 Vss 0.00213842f
c123 63 Vss 0.00546856f
c124 59 Vss 0.00725053f
c125 54 Vss 0.00546856f
c126 45 Vss 1.15207e-19
c127 43 Vss 0.0351228f
c128 42 Vss 0.100955f
c129 33 Vss 0.035919f
c130 32 Vss 0.100953f
c131 14 Vss 0.00143442f
c132 9 Vss 0.266831f
c133 5 Vss 0.270069f
r134 98 103 0.326018
r135 97 98 4.58464
r136 93 97 0.655813
r137 93 95 1.82344
r138 92 101 0.494161
r139 91 103 0.326018
r140 91 92 13.0037
r141 87 101 0.128424
r142 87 89 5.2515
r143 85 114 1.16709
r144 83 85 2.16729
r145 82 100 0.494161
r146 81 101 0.494161
r147 81 82 7.46046
r148 79 109 1.16709
r149 77 100 0.128424
r150 77 79 2.16729
r151 75 100 0.494161
r152 75 76 4.37625
r153 71 99 0.0828784
r154 71 73 1.82344
r155 69 83 0.652036
r156 69 70 10.1279
r157 68 76 0.652036
r158 67 99 0.551426
r159 67 68 14.7125
r160 66 99 0.551426
r161 65 70 0.652036
r162 65 66 4.58464
r163 63 95 1.16709
r164 59 89 1.16709
r165 54 73 1.16709
r166 45 114 0.0476429
r167 43 45 1.45875
r168 42 46 0.652036
r169 42 45 1.45875
r170 39 43 0.652036
r171 35 109 0.0476429
r172 33 35 1.45875
r173 32 36 0.652036
r174 32 35 1.45875
r175 29 33 0.652036
r176 16 63 0.185659
r177 14 59 0.185659
r178 12 59 0.185659
r179 9 46 3.8511
r180 9 39 3.8511
r181 5 36 3.8511
r182 5 29 3.8511
r183 2 54 0.185659
.ends

.subckt PM_G4_XNOR2_N2_VSS 3 6 8 11 14 16 32 33 42 43 54 59 63 66 71 76 81 87 96
+ 101 114 116 117 118 123 124 129 137 142 143 144 146 Vss
c87 144 Vss 3.75522e-19
c88 143 Vss 4.28045e-19
c89 142 Vss 0.00380395f
c90 137 Vss 0.00119929f
c91 129 Vss 0.0129925f
c92 124 Vss 8.20954e-19
c93 123 Vss 0.00416713f
c94 118 Vss 8.42922e-19
c95 117 Vss 0.00171404f
c96 116 Vss 0.00154361f
c97 114 Vss 0.00516329f
c98 101 Vss 0.00400427f
c99 96 Vss 0.00412244f
c100 87 Vss 1.41859e-19
c101 81 Vss 0.00270839f
c102 76 Vss 8.07404e-19
c103 71 Vss 0.00125472f
c104 66 Vss 0.00178947f
c105 63 Vss 0.00389308f
c106 59 Vss 0.00728678f
c107 54 Vss 0.0039211f
c108 43 Vss 0.0342891f
c109 42 Vss 0.100066f
c110 35 Vss 1.95386e-19
c111 33 Vss 0.0350852f
c112 32 Vss 0.0990713f
c113 14 Vss 0.00143442f
c114 11 Vss 0.269838f
c115 3 Vss 0.266926f
r116 142 146 0.349767
r117 141 142 4.58464
r118 137 146 0.306046
r119 130 144 0.494161
r120 129 141 0.652036
r121 125 144 0.128424
r122 123 133 0.652036
r123 123 124 10.1279
r124 119 143 0.0828784
r125 117 144 0.494161
r126 117 118 4.37625
r127 116 124 0.652036
r128 115 143 0.551426
r129 115 116 4.58464
r130 114 143 0.551426
r131 113 118 0.652036
r132 113 114 14.7125
r133 87 137 1.82344
r134 81 129 13.5872
r135 81 130 8.04396
r136 81 84 5.79332
r137 76 101 1.16709
r138 76 133 2.16729
r139 71 96 1.16709
r140 71 125 2.16729
r141 66 119 1.82344
r142 63 87 1.16709
r143 59 84 1.16709
r144 54 66 1.16709
r145 45 101 0.0476429
r146 43 45 1.45875
r147 42 46 0.652036
r148 42 45 1.45875
r149 39 43 0.652036
r150 35 96 0.0476429
r151 33 35 1.45875
r152 32 36 0.652036
r153 32 35 1.45875
r154 29 33 0.652036
r155 16 63 0.185659
r156 14 59 0.185659
r157 11 46 3.8511
r158 11 39 3.8511
r159 8 59 0.185659
r160 6 54 0.185659
r161 3 36 3.8511
r162 3 29 3.8511
.ends

.subckt PM_G4_XNOR2_N2_A 2 4 7 10 21 24 28 39 48 53 56 61 66 71 76 84 Vss
c57 84 Vss 4.74028e-19
c58 76 Vss 8.09766e-19
c59 71 Vss 0.00526551f
c60 66 Vss 0.00379683f
c61 61 Vss 0.00265207f
c62 56 Vss 0.0049943f
c63 53 Vss 8.5599e-19
c64 48 Vss 0.126052f
c65 43 Vss 0.0296526f
c66 39 Vss 1.95944e-19
c67 28 Vss 0.152877f
c68 24 Vss 1.05421e-19
c69 21 Vss 0.169632f
c70 18 Vss 0.12596f
c71 16 Vss 0.0247918f
c72 10 Vss 0.121972f
c73 7 Vss 0.324361f
c74 4 Vss 0.138512f
r75 80 84 0.652036
r76 61 76 1.16709
r77 61 84 5.20982
r78 56 71 1.16709
r79 56 80 9.54439
r80 53 66 1.16709
r81 47 71 0.0238214
r82 47 48 2.334
r83 44 47 2.20433
r84 39 76 0.404964
r85 33 48 0.00605528
r86 31 44 0.00605528
r87 29 43 0.494161
r88 28 30 0.652036
r89 28 29 4.84305
r90 25 43 0.128424
r91 24 66 0.0476429
r92 22 24 0.326018
r93 22 24 0.1167
r94 21 43 0.494161
r95 21 24 6.7686
r96 18 66 0.357321
r97 16 24 0.326018
r98 16 18 0.40845
r99 10 39 3.32595
r100 7 33 3.8511
r101 7 31 3.8511
r102 7 30 3.8511
r103 4 25 3.8511
r104 2 18 3.44265
.ends

.subckt PM_G4_XNOR2_N2_NET1 2 4 7 10 30 31 35 41 44 49 58 66 Vss
c34 66 Vss 2.19199e-19
c35 58 Vss 0.0058571f
c36 49 Vss 0.00612925f
c37 44 Vss 0.00128347f
c38 41 Vss 0.00534332f
c39 35 Vss 0.103384f
c40 31 Vss 0.12896f
c41 30 Vss 1.02017e-19
c42 10 Vss 0.236304f
c43 7 Vss 0.381296f
c44 4 Vss 0.00143442f
r45 62 66 0.652036
r46 49 58 1.16709
r47 49 66 13.8373
r48 44 62 2.50071
r49 41 44 1.16709
r50 33 35 1.70187
r51 30 58 0.0238214
r52 30 31 2.20433
r53 27 30 2.334
r54 25 35 0.17282
r55 24 31 0.00605528
r56 21 33 0.17282
r57 18 27 0.00605528
r58 10 21 7.06035
r59 7 25 5.7183
r60 7 24 3.8511
r61 7 18 3.8511
r62 4 41 0.185659
r63 2 41 0.185659
.ends

.subckt PM_G4_XNOR2_N2_NET3 2 4 6 9 21 22 33 39 42 47 56 74 Vss
c49 74 Vss 3.4517e-19
c50 56 Vss 0.0039047f
c51 47 Vss 0.00714759f
c52 42 Vss 0.00198779f
c53 39 Vss 0.00534332f
c54 33 Vss 0.12548f
c55 22 Vss 0.0340569f
c56 21 Vss 0.175814f
c57 9 Vss 0.464757f
c58 6 Vss 0.145805f
c59 4 Vss 0.00143442f
r60 70 74 0.655813
r61 47 56 1.16709
r62 47 74 12.0712
r63 42 70 2.41736
r64 39 42 1.16709
r65 32 56 0.0238214
r66 32 33 2.26917
r67 29 32 2.26917
r68 26 33 0.00605528
r69 24 29 0.00605528
r70 21 23 0.652036
r71 21 22 4.84305
r72 18 22 0.652036
r73 9 26 3.8511
r74 9 24 3.8511
r75 9 23 8.7525
r76 6 18 4.25955
r77 4 39 0.185659
r78 2 39 0.185659
.ends

.subckt PM_G4_XNOR2_N2_B 2 4 7 10 19 20 28 31 33 37 38 48 52 58 61 Vss
c36 61 Vss 0.0281739f
c37 58 Vss 0.00110612f
c38 52 Vss 0.136411f
c39 48 Vss 0.0595342f
c40 38 Vss 0.0333783f
c41 37 Vss 0.090268f
c42 33 Vss 0.0442143f
c43 31 Vss 9.80304e-20
c44 28 Vss 0.0899896f
c45 20 Vss 0.0348277f
c46 19 Vss 0.169632f
c47 10 Vss 0.209756f
c48 7 Vss 0.322768f
c49 4 Vss 0.125964f
c50 2 Vss 0.138383f
r51 55 61 1.16709
r52 55 58 0.0729375
r53 50 52 4.53833
r54 47 48 1.167
r55 42 52 0.00605528
r56 37 39 0.652036
r57 37 38 2.04225
r58 35 48 0.0685365
r59 34 50 0.00605528
r60 33 38 0.652036
r61 32 47 0.0685365
r62 32 33 1.69215
r63 31 61 0.181909
r64 29 61 0.494161
r65 29 31 0.1167
r66 28 47 0.5835
r67 28 31 3.55935
r68 23 61 0.128424
r69 23 61 0.40845
r70 22 61 0.181909
r71 20 22 6.7686
r72 19 61 0.494161
r73 19 22 0.1167
r74 16 20 0.652036
r75 10 39 6.3018
r76 7 42 3.8511
r77 7 35 3.8511
r78 7 34 3.8511
r79 4 61 3.44265
r80 2 16 3.8511
.ends

.subckt PM_G4_XNOR2_N2_Z 2 4 6 8 23 27 30 33 Vss
c29 30 Vss 0.00338645f
c30 27 Vss 0.0063256f
c31 23 Vss 0.00620875f
c32 8 Vss 0.00143442f
c33 6 Vss 0.00143442f
r34 33 35 4.668
r35 30 33 5.45989
r36 27 35 1.16709
r37 23 30 1.16709
r38 8 27 0.185659
r39 6 23 0.185659
r40 4 27 0.185659
r41 2 23 0.185659
.ends

.subckt G4_XNOR2_N2  VDD VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI16.X0 N_NET1_XI16.X0_D N_VSS_XI16.X0_PGD N_B_XI16.X0_CG N_VSS_XI16.X0_PGD
+ N_VDD_XI16.X0_S TIGFET_HPNW8
XI12.X0 N_NET3_XI12.X0_D N_VDD_XI12.X0_PGD N_A_XI12.X0_CG N_VDD_XI12.X0_PGD
+ N_VSS_XI12.X0_S TIGFET_HPNW8
XI18.X0 N_NET1_XI18.X0_D N_VDD_XI18.X0_PGD N_B_XI18.X0_CG N_VDD_XI18.X0_PGD
+ N_VSS_XI18.X0_S TIGFET_HPNW8
XI13.X0 N_NET3_XI13.X0_D N_VSS_XI13.X0_PGD N_A_XI13.X0_CG N_VSS_XI13.X0_PGD
+ N_VDD_XI13.X0_S TIGFET_HPNW8
XI17.X0 N_Z_XI17.X0_D N_B_XI17.X0_PGD N_NET3_XI17.X0_CG N_B_XI17.X0_PGD
+ N_VSS_XI17.X0_S TIGFET_HPNW8
XI14.X0 N_Z_XI14.X0_D N_A_XI14.X0_PGD N_B_XI14.X0_CG N_A_XI14.X0_PGD
+ N_VDD_XI14.X0_S TIGFET_HPNW8
XI19.X0 N_Z_XI19.X0_D N_NET1_XI19.X0_PGD N_A_XI19.X0_CG N_NET1_XI19.X0_PGD
+ N_VSS_XI19.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_NET3_XI15.X0_PGD N_NET1_XI15.X0_CG N_NET3_XI15.X0_PGD
+ N_VDD_XI15.X0_S TIGFET_HPNW8
*
x_PM_G4_XNOR2_N2_VDD N_VDD_XI16.X0_S N_VDD_XI12.X0_PGD N_VDD_XI18.X0_PGD
+ N_VDD_XI13.X0_S N_VDD_XI14.X0_S N_VDD_XI15.X0_S N_VDD_c_9_p N_VDD_c_23_p
+ N_VDD_c_5_p N_VDD_c_89_p N_VDD_c_65_p N_VDD_c_11_p N_VDD_c_96_p N_VDD_c_7_p
+ N_VDD_c_12_p N_VDD_c_6_p N_VDD_c_40_p N_VDD_c_13_p N_VDD_c_14_p N_VDD_c_44_p
+ N_VDD_c_19_p N_VDD_c_10_p N_VDD_c_17_p N_VDD_c_4_p N_VDD_c_54_p N_VDD_c_27_p
+ N_VDD_c_72_p N_VDD_c_37_p N_VDD_c_43_p VDD N_VDD_c_22_p N_VDD_c_18_p Vss
+ PM_G4_XNOR2_N2_VDD
x_PM_G4_XNOR2_N2_VSS N_VSS_XI16.X0_PGD N_VSS_XI12.X0_S N_VSS_XI18.X0_S
+ N_VSS_XI13.X0_PGD N_VSS_XI17.X0_S N_VSS_XI19.X0_S N_VSS_c_109_n N_VSS_c_111_n
+ N_VSS_c_157_p N_VSS_c_113_n N_VSS_c_173_p N_VSS_c_115_n N_VSS_c_185_p
+ N_VSS_c_116_n N_VSS_c_119_n N_VSS_c_123_n N_VSS_c_127_n N_VSS_c_131_n
+ N_VSS_c_132_n N_VSS_c_136_n N_VSS_c_139_n N_VSS_c_142_n N_VSS_c_143_n
+ N_VSS_c_144_n N_VSS_c_145_n N_VSS_c_148_n N_VSS_c_149_n N_VSS_c_150_n
+ N_VSS_c_169_p N_VSS_c_151_n N_VSS_c_152_n VSS Vss PM_G4_XNOR2_N2_VSS
x_PM_G4_XNOR2_N2_A N_A_XI12.X0_CG N_A_XI13.X0_CG N_A_XI14.X0_PGD N_A_XI19.X0_CG
+ N_A_c_193_n N_A_c_195_n N_A_c_196_n N_A_c_220_p N_A_c_197_n A N_A_c_201_n
+ N_A_c_221_p N_A_c_203_n N_A_c_206_n N_A_c_219_p N_A_c_217_n Vss
+ PM_G4_XNOR2_N2_A
x_PM_G4_XNOR2_N2_NET1 N_NET1_XI16.X0_D N_NET1_XI18.X0_D N_NET1_XI19.X0_PGD
+ N_NET1_XI15.X0_CG N_NET1_c_268_n N_NET1_c_281_p N_NET1_c_274_p N_NET1_c_249_n
+ N_NET1_c_252_n N_NET1_c_255_n N_NET1_c_271_n N_NET1_c_263_n Vss
+ PM_G4_XNOR2_N2_NET1
x_PM_G4_XNOR2_N2_NET3 N_NET3_XI12.X0_D N_NET3_XI13.X0_D N_NET3_XI17.X0_CG
+ N_NET3_XI15.X0_PGD N_NET3_c_306_n N_NET3_c_323_p N_NET3_c_284_n N_NET3_c_285_n
+ N_NET3_c_286_n N_NET3_c_289_n N_NET3_c_292_n N_NET3_c_294_n Vss
+ PM_G4_XNOR2_N2_NET3
x_PM_G4_XNOR2_N2_B N_B_XI16.X0_CG N_B_XI18.X0_CG N_B_XI17.X0_PGD N_B_XI14.X0_CG
+ N_B_c_334_n N_B_c_349_n N_B_c_336_n N_B_c_337_n N_B_c_361_n N_B_c_357_n
+ N_B_c_351_n N_B_c_365_n N_B_c_338_n B N_B_c_341_n Vss PM_G4_XNOR2_N2_B
x_PM_G4_XNOR2_N2_Z N_Z_XI17.X0_D N_Z_XI14.X0_D N_Z_XI19.X0_D N_Z_XI15.X0_D
+ N_Z_c_378_n N_Z_c_368_n N_Z_c_373_n Z Vss PM_G4_XNOR2_N2_Z
cc_1 N_VDD_XI12.X0_PGD N_VSS_XI16.X0_PGD 2.89249e-19
cc_2 N_VDD_XI18.X0_PGD N_VSS_XI16.X0_PGD 0.00196286f
cc_3 N_VDD_XI12.X0_PGD N_VSS_XI13.X0_PGD 0.0019593f
cc_4 N_VDD_c_4_p N_VSS_XI13.X0_PGD 2.22629e-19
cc_5 N_VDD_c_5_p N_VSS_c_109_n 0.00196286f
cc_6 N_VDD_c_6_p N_VSS_c_109_n 3.9313e-19
cc_7 N_VDD_c_7_p N_VSS_c_111_n 2.76462e-19
cc_8 N_VDD_c_6_p N_VSS_c_111_n 3.9313e-19
cc_9 N_VDD_c_9_p N_VSS_c_113_n 0.0019593f
cc_10 N_VDD_c_10_p N_VSS_c_113_n 3.9313e-19
cc_11 N_VDD_c_11_p N_VSS_c_115_n 3.13688e-19
cc_12 N_VDD_c_12_p N_VSS_c_116_n 0.00187494f
cc_13 N_VDD_c_13_p N_VSS_c_116_n 5.06564e-19
cc_14 N_VDD_c_14_p N_VSS_c_116_n 4.5625e-19
cc_15 N_VDD_c_7_p N_VSS_c_119_n 4.35319e-19
cc_16 N_VDD_c_6_p N_VSS_c_119_n 0.00141228f
cc_17 N_VDD_c_17_p N_VSS_c_119_n 8.69067e-19
cc_18 N_VDD_c_18_p N_VSS_c_119_n 3.48267e-19
cc_19 N_VDD_c_19_p N_VSS_c_123_n 9.53862e-19
cc_20 N_VDD_c_10_p N_VSS_c_123_n 0.00161703f
cc_21 N_VDD_c_4_p N_VSS_c_123_n 0.00227772f
cc_22 N_VDD_c_22_p N_VSS_c_123_n 3.48267e-19
cc_23 N_VDD_c_23_p N_VSS_c_127_n 2.38046e-19
cc_24 N_VDD_c_6_p N_VSS_c_127_n 0.00534412f
cc_25 N_VDD_c_4_p N_VSS_c_127_n 3.34043e-19
cc_26 N_VDD_c_18_p N_VSS_c_127_n 9.58524e-19
cc_27 N_VDD_c_27_p N_VSS_c_131_n 2.11881e-19
cc_28 N_VDD_c_7_p N_VSS_c_132_n 3.66936e-19
cc_29 N_VDD_c_6_p N_VSS_c_132_n 0.00114511f
cc_30 N_VDD_c_17_p N_VSS_c_132_n 3.99794e-19
cc_31 N_VDD_c_18_p N_VSS_c_132_n 6.489e-19
cc_32 N_VDD_c_10_p N_VSS_c_136_n 2.26455e-19
cc_33 N_VDD_c_4_p N_VSS_c_136_n 9.55322e-19
cc_34 N_VDD_c_22_p N_VSS_c_136_n 6.46219e-19
cc_35 N_VDD_c_7_p N_VSS_c_139_n 0.00309754f
cc_36 N_VDD_c_12_p N_VSS_c_139_n 0.00766101f
cc_37 N_VDD_c_37_p N_VSS_c_139_n 0.0010706f
cc_38 N_VDD_c_12_p N_VSS_c_142_n 0.0033176f
cc_39 N_VDD_c_6_p N_VSS_c_143_n 0.00345383f
cc_40 N_VDD_c_40_p N_VSS_c_144_n 0.00107685f
cc_41 N_VDD_c_14_p N_VSS_c_145_n 0.0035394f
cc_42 N_VDD_c_10_p N_VSS_c_145_n 0.00604286f
cc_43 N_VDD_c_43_p N_VSS_c_145_n 0.00103916f
cc_44 N_VDD_c_44_p N_VSS_c_148_n 0.0010609f
cc_45 N_VDD_c_6_p N_VSS_c_149_n 0.00459995f
cc_46 N_VDD_c_27_p N_VSS_c_150_n 0.00107435f
cc_47 N_VDD_c_12_p N_VSS_c_151_n 9.16632e-19
cc_48 N_VDD_c_6_p N_VSS_c_152_n 7.74609e-19
cc_49 N_VDD_c_4_p N_A_XI14.X0_PGD 2.06119e-19
cc_50 N_VDD_XI12.X0_PGD N_A_c_193_n 4.07423e-19
cc_51 N_VDD_XI18.X0_PGD N_A_c_193_n 2.2186e-19
cc_52 N_VDD_c_22_p N_A_c_195_n 9.45508e-19
cc_53 N_VDD_XI18.X0_PGD N_A_c_196_n 2.2186e-19
cc_54 N_VDD_c_54_p N_A_c_197_n 6.28504e-19
cc_55 N_VDD_c_12_p A 5.04211e-19
cc_56 N_VDD_c_19_p A 4.35492e-19
cc_57 N_VDD_c_22_p A 3.2351e-19
cc_58 N_VDD_c_4_p N_A_c_201_n 0.00256103f
cc_59 N_VDD_c_54_p N_A_c_201_n 0.00191796f
cc_60 N_VDD_c_12_p N_A_c_203_n 6.26183e-19
cc_61 N_VDD_c_19_p N_A_c_203_n 3.43988e-19
cc_62 N_VDD_c_22_p N_A_c_203_n 2.68747e-19
cc_63 N_VDD_c_4_p N_A_c_206_n 9.84209e-19
cc_64 N_VDD_c_54_p N_A_c_206_n 2.68554e-19
cc_65 N_VDD_c_65_p N_NET1_c_249_n 3.43419e-19
cc_66 N_VDD_c_6_p N_NET1_c_249_n 3.4118e-19
cc_67 N_VDD_c_13_p N_NET1_c_249_n 3.72199e-19
cc_68 N_VDD_c_65_p N_NET1_c_252_n 3.48267e-19
cc_69 N_VDD_c_6_p N_NET1_c_252_n 3.98099e-19
cc_70 N_VDD_c_13_p N_NET1_c_252_n 5.226e-19
cc_71 N_VDD_c_17_p N_NET1_c_255_n 0.00115819f
cc_72 N_VDD_c_72_p N_NET3_XI15.X0_PGD 2.91063e-19
cc_73 N_VDD_c_54_p N_NET3_c_284_n 8.60495e-19
cc_74 N_VDD_c_11_p N_NET3_c_285_n 3.43419e-19
cc_75 N_VDD_c_11_p N_NET3_c_286_n 3.48267e-19
cc_76 N_VDD_c_10_p N_NET3_c_286_n 4.34701e-19
cc_77 N_VDD_c_4_p N_NET3_c_286_n 0.00100809f
cc_78 N_VDD_c_4_p N_NET3_c_289_n 0.00119634f
cc_79 N_VDD_c_54_p N_NET3_c_289_n 0.00298078f
cc_80 N_VDD_c_72_p N_NET3_c_289_n 7.77543e-19
cc_81 N_VDD_c_54_p N_NET3_c_292_n 0.00118178f
cc_82 N_VDD_c_72_p N_NET3_c_292_n 3.66936e-19
cc_83 N_VDD_c_19_p N_NET3_c_294_n 2.94103e-19
cc_84 N_VDD_c_12_p N_B_XI16.X0_CG 2.61808e-19
cc_85 N_VDD_XI18.X0_PGD N_B_XI17.X0_PGD 0.00190378f
cc_86 N_VDD_XI12.X0_PGD N_B_c_334_n 2.2186e-19
cc_87 N_VDD_XI18.X0_PGD N_B_c_334_n 4.07423e-19
cc_88 N_VDD_XI18.X0_PGD N_B_c_336_n 4.08222e-19
cc_89 N_VDD_c_89_p N_B_c_337_n 9.08628e-19
cc_90 N_VDD_c_23_p N_B_c_338_n 0.00168656f
cc_91 N_VDD_c_17_p B 3.02102e-19
cc_92 N_VDD_c_18_p B 3.2351e-19
cc_93 N_VDD_c_17_p N_B_c_341_n 3.36818e-19
cc_94 N_VDD_c_18_p N_B_c_341_n 2.68747e-19
cc_95 N_VDD_c_11_p N_Z_c_368_n 3.43419e-19
cc_96 N_VDD_c_96_p N_Z_c_368_n 3.43419e-19
cc_97 N_VDD_c_4_p N_Z_c_368_n 3.48267e-19
cc_98 N_VDD_c_54_p N_Z_c_368_n 3.4118e-19
cc_99 N_VDD_c_27_p N_Z_c_368_n 3.72199e-19
cc_100 N_VDD_c_11_p N_Z_c_373_n 3.48267e-19
cc_101 N_VDD_c_96_p N_Z_c_373_n 3.48267e-19
cc_102 N_VDD_c_4_p N_Z_c_373_n 4.85404e-19
cc_103 N_VDD_c_54_p N_Z_c_373_n 5.96492e-19
cc_104 N_VDD_c_27_p N_Z_c_373_n 8.21216e-19
cc_105 N_VSS_XI13.X0_PGD N_A_XI14.X0_PGD 0.00164979f
cc_106 N_VSS_XI16.X0_PGD N_A_c_193_n 2.2186e-19
cc_107 N_VSS_XI13.X0_PGD N_A_c_193_n 4.04227e-19
cc_108 N_VSS_XI13.X0_PGD N_A_c_196_n 4.08222e-19
cc_109 N_VSS_c_157_p N_A_c_197_n 0.00164979f
cc_110 N_VSS_c_123_n N_A_c_201_n 3.87149e-19
cc_111 N_VSS_c_139_n N_A_c_201_n 4.99859e-19
cc_112 N_VSS_c_132_n N_A_c_203_n 2.38312e-19
cc_113 N_VSS_c_136_n N_A_c_206_n 6.52904e-19
cc_114 N_VSS_c_149_n N_A_c_217_n 6.07247e-19
cc_115 N_VSS_c_115_n N_NET1_c_249_n 3.43419e-19
cc_116 N_VSS_c_127_n N_NET1_c_249_n 3.48267e-19
cc_117 N_VSS_c_115_n N_NET1_c_252_n 3.48267e-19
cc_118 N_VSS_c_127_n N_NET1_c_252_n 0.00138658f
cc_119 N_VSS_c_127_n N_NET1_c_255_n 0.00157945f
cc_120 N_VSS_c_149_n N_NET1_c_255_n 0.0182344f
cc_121 N_VSS_c_169_p N_NET1_c_255_n 0.0011475f
cc_122 N_VSS_c_119_n N_NET1_c_263_n 0.00193107f
cc_123 N_VSS_c_139_n N_NET1_c_263_n 0.00107322f
cc_124 N_VSS_c_149_n N_NET1_c_263_n 0.00164616f
cc_125 N_VSS_c_173_p N_NET3_c_285_n 3.43419e-19
cc_126 N_VSS_c_173_p N_NET3_c_286_n 3.48267e-19
cc_127 N_VSS_c_116_n N_NET3_c_286_n 0.0011211f
cc_128 N_VSS_c_142_n N_NET3_c_286_n 4.15771e-19
cc_129 N_VSS_c_145_n N_NET3_c_286_n 2.79692e-19
cc_130 N_VSS_c_123_n N_NET3_c_289_n 0.00136387f
cc_131 N_VSS_c_145_n N_NET3_c_294_n 4.73555e-19
cc_132 N_VSS_XI16.X0_PGD N_B_c_334_n 4.04227e-19
cc_133 N_VSS_XI13.X0_PGD N_B_c_334_n 2.2186e-19
cc_134 N_VSS_XI13.X0_PGD N_B_c_336_n 2.2186e-19
cc_135 N_VSS_c_127_n N_B_c_338_n 2.49315e-19
cc_136 N_VSS_c_115_n N_Z_c_378_n 3.43419e-19
cc_137 N_VSS_c_185_p N_Z_c_378_n 3.43419e-19
cc_138 N_VSS_c_127_n N_Z_c_378_n 3.48267e-19
cc_139 N_VSS_c_131_n N_Z_c_378_n 3.48267e-19
cc_140 N_VSS_c_115_n N_Z_c_373_n 3.48267e-19
cc_141 N_VSS_c_185_p N_Z_c_373_n 3.48267e-19
cc_142 N_VSS_c_127_n N_Z_c_373_n 8.69457e-19
cc_143 N_VSS_c_131_n N_Z_c_373_n 5.71987e-19
cc_144 N_A_XI19.X0_CG N_NET1_XI19.X0_PGD 5.00154e-19
cc_145 N_A_c_219_p N_NET1_XI19.X0_PGD 0.00253213f
cc_146 N_A_c_220_p N_NET1_c_268_n 9.11431e-19
cc_147 N_A_c_221_p N_NET1_c_255_n 0.00300988f
cc_148 N_A_c_217_n N_NET1_c_255_n 8.60245e-19
cc_149 N_A_c_221_p N_NET1_c_271_n 3.14782e-19
cc_150 N_A_c_219_p N_NET1_c_271_n 2.68747e-19
cc_151 N_A_c_219_p N_NET3_XI17.X0_CG 2.16281e-19
cc_152 N_A_XI14.X0_PGD N_NET3_XI15.X0_PGD 0.00174198f
cc_153 N_A_c_196_n N_NET3_XI15.X0_PGD 3.14428e-19
cc_154 N_A_c_219_p N_NET3_XI15.X0_PGD 4.34237e-19
cc_155 N_A_XI14.X0_PGD N_NET3_c_306_n 4.63684e-19
cc_156 N_A_c_197_n N_NET3_c_284_n 0.00174198f
cc_157 N_A_c_193_n N_NET3_c_285_n 6.32063e-19
cc_158 N_A_c_201_n N_NET3_c_286_n 9.99037e-19
cc_159 N_A_c_201_n N_NET3_c_289_n 0.00251926f
cc_160 N_A_c_221_p N_NET3_c_289_n 0.00147102f
cc_161 N_A_c_206_n N_NET3_c_289_n 3.44698e-19
cc_162 N_A_c_220_p N_NET3_c_292_n 4.02896e-19
cc_163 N_A_c_201_n N_NET3_c_292_n 3.44698e-19
cc_164 N_A_c_206_n N_NET3_c_292_n 6.70706e-19
cc_165 N_A_c_196_n N_B_XI14.X0_CG 0.003858f
cc_166 N_A_c_193_n N_B_c_334_n 0.00500727f
cc_167 N_A_c_203_n N_B_c_349_n 6.36314e-19
cc_168 N_A_c_196_n N_B_c_336_n 0.00268264f
cc_169 N_A_c_196_n N_B_c_351_n 0.00354125f
cc_170 N_A_c_217_n B 2.16641e-19
cc_171 N_A_c_193_n N_B_c_341_n 0.00152783f
cc_172 N_A_c_201_n N_Z_c_373_n 0.00406991f
cc_173 N_A_c_221_p N_Z_c_373_n 0.00267623f
cc_174 N_A_c_219_p N_Z_c_373_n 0.00100289f
cc_175 N_NET1_XI19.X0_PGD N_NET3_XI17.X0_CG 3.24817e-19
cc_176 N_NET1_c_274_p N_NET3_XI15.X0_PGD 0.00863799f
cc_177 N_NET1_XI19.X0_PGD N_NET3_c_306_n 0.00333245f
cc_178 N_NET1_c_249_n N_NET3_c_285_n 2.31842e-19
cc_179 N_NET1_XI19.X0_PGD N_B_XI17.X0_PGD 0.00216194f
cc_180 N_NET1_XI15.X0_CG N_B_XI14.X0_CG 2.72501e-19
cc_181 N_NET1_c_249_n N_B_c_334_n 6.32063e-19
cc_182 N_NET1_c_274_p N_B_c_357_n 2.72501e-19
cc_183 N_NET1_c_281_p N_B_c_338_n 0.00193608f
cc_184 N_NET1_c_255_n N_Z_c_373_n 3.07539e-19
cc_185 N_NET3_XI17.X0_CG N_B_XI17.X0_PGD 0.00201028f
cc_186 N_NET3_c_306_n N_B_XI17.X0_PGD 0.00163252f
cc_187 N_NET3_XI15.X0_PGD N_B_c_361_n 3.23792e-19
cc_188 N_NET3_c_323_p N_B_c_361_n 5.75886e-19
cc_189 N_NET3_XI15.X0_PGD N_B_c_357_n 0.00310335f
cc_190 N_NET3_c_323_p N_B_c_357_n 0.00192667f
cc_191 N_NET3_c_323_p N_B_c_365_n 0.00201028f
cc_192 N_NET3_c_306_n N_Z_c_378_n 6.54859e-19
cc_193 N_NET3_c_306_n N_Z_c_368_n 2.54846e-19
cc_194 N_NET3_XI15.X0_PGD N_Z_c_373_n 0.00129454f
cc_195 N_NET3_c_306_n N_Z_c_373_n 2.46041e-19
cc_196 N_NET3_c_289_n N_Z_c_373_n 2.36895e-19
cc_197 N_B_c_357_n N_Z_c_373_n 9.47639e-19
cc_198 B N_Z_c_373_n 2.02757e-19
*
.ends
*
*
.subckt XNOR2_HPNW8 A B Y VDD VSS
xgate (VDD VSS A B Y) G4_XNOR2_N2
.ends
*
* File: G5_XNOR3_N2.pex.netlist
* Created: Mon Mar 28 15:31:24 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XNOR3_N2_VDD 2 3 5 8 10 11 29 30 41 42 44 53 54 65 69 74 83 85 86
+ 87 90 92 96 99 102 104 108 110 114 118 120 122 124 125 131 140 145 Vss
c116 145 Vss 0.00470693f
c117 140 Vss 0.00487376f
c118 131 Vss 0.00472091f
c119 125 Vss 2.39889e-19
c120 124 Vss 4.91772e-19
c121 123 Vss 5.21614e-19
c122 120 Vss 4.52364e-19
c123 118 Vss 0.00162316f
c124 114 Vss 4.81041e-19
c125 110 Vss 0.00631991f
c126 108 Vss 9.42823e-19
c127 104 Vss 0.00578311f
c128 102 Vss 0.00174133f
c129 99 Vss 0.00271006f
c130 96 Vss 0.00486611f
c131 92 Vss 0.00657264f
c132 90 Vss 0.00151669f
c133 87 Vss 8.67714e-19
c134 86 Vss 0.0090076f
c135 85 Vss 0.0105886f
c136 83 Vss 0.00212071f
c137 74 Vss 0.00377995f
c138 69 Vss 0.0039448f
c139 65 Vss 0.00373195f
c140 54 Vss 0.035607f
c141 53 Vss 0.100823f
c142 44 Vss 8.7772e-20
c143 42 Vss 0.0356105f
c144 41 Vss 0.101295f
c145 30 Vss 0.0346327f
c146 29 Vss 0.0990915f
c147 11 Vss 0.269218f
c148 5 Vss 0.27009f
c149 3 Vss 0.232895f
r150 116 118 5.2515
r151 114 145 1.16709
r152 112 114 2.16729
r153 111 125 0.494161
r154 110 116 0.652036
r155 110 111 7.46046
r156 108 140 1.16709
r157 106 125 0.128424
r158 106 108 2.16729
r159 105 124 0.494161
r160 104 112 0.652036
r161 104 105 10.3363
r162 100 123 0.0828784
r163 100 102 2.00578
r164 99 124 0.128424
r165 98 123 0.551426
r166 98 99 4.58464
r167 96 131 1.16709
r168 94 123 0.551426
r169 94 96 7.25207
r170 93 122 0.326018
r171 92 124 0.494161
r172 92 93 10.1279
r173 88 120 0.0828784
r174 88 90 1.82344
r175 86 125 0.494161
r176 86 87 15.8795
r177 85 122 0.326018
r178 84 120 0.551426
r179 84 85 15.5878
r180 83 120 0.551426
r181 82 87 0.652036
r182 82 83 4.58464
r183 74 118 1.16709
r184 69 102 1.16709
r185 65 90 1.16709
r186 56 145 0.0476429
r187 54 56 1.45875
r188 53 57 0.652036
r189 53 56 1.45875
r190 49 54 0.652036
r191 44 140 0.0476429
r192 42 44 1.45875
r193 41 45 0.652036
r194 41 44 1.45875
r195 37 42 0.652036
r196 32 131 0.238214
r197 30 32 1.45875
r198 29 33 0.652036
r199 29 32 1.45875
r200 25 30 0.652036
r201 11 57 3.8511
r202 11 49 3.8511
r203 10 74 0.185659
r204 8 69 0.185659
r205 5 45 3.8511
r206 5 37 3.8511
r207 3 33 3.1509
r208 3 25 3.1509
r209 2 65 0.185659
.ends

.subckt PM_G5_XNOR3_N2_C 2 4 6 8 20 23 32 40 43 47 52 57 67 86 94 100 Vss
c51 100 Vss 3.07518e-19
c52 94 Vss 0.00534351f
c53 86 Vss 0.010496f
c54 67 Vss 0.00399096f
c55 57 Vss 0.00459151f
c56 52 Vss 0.00198824f
c57 47 Vss 0.00148308f
c58 43 Vss 0.00113252f
c59 32 Vss 0.00492048f
c60 23 Vss 9.8832e-20
c61 20 Vss 0.221837f
c62 17 Vss 0.126125f
c63 15 Vss 0.0247918f
c64 4 Vss 0.133869f
r65 95 100 0.494161
r66 94 96 0.652036
r67 94 95 10.3363
r68 90 100 0.128424
r69 86 100 0.494161
r70 57 60 0.05
r71 52 67 1.16709
r72 52 96 2.37568
r73 47 90 2.45904
r74 43 60 1.16709
r75 43 86 25.2989
r76 40 43 0.0364688
r77 37 67 0.1
r78 32 47 1.16709
r79 23 57 0.0476429
r80 21 23 0.326018
r81 21 23 0.1167
r82 20 24 0.652036
r83 20 23 6.7686
r84 17 57 0.357321
r85 15 23 0.326018
r86 15 17 0.40845
r87 8 37 0.185659
r88 6 32 0.185659
r89 4 24 3.8511
r90 2 17 3.44265
.ends

.subckt PM_G5_XNOR3_N2_VSS 1 4 6 7 9 12 29 32 41 42 53 54 56 66 70 79 84 89 94
+ 99 102 105 114 119 128 130 131 132 137 138 143 151 159 160 161 Vss
c126 161 Vss 3.75522e-19
c127 160 Vss 3.88979e-19
c128 159 Vss 4.4306e-19
c129 143 Vss 0.00346584f
c130 138 Vss 8.41415e-19
c131 137 Vss 0.00629302f
c132 132 Vss 8.38477e-19
c133 131 Vss 0.00556756f
c134 130 Vss 0.00421531f
c135 128 Vss 0.00274186f
c136 119 Vss 0.00392167f
c137 114 Vss 0.00408379f
c138 105 Vss 0.00489622f
c139 102 Vss 0.00348146f
c140 99 Vss 0.00311148f
c141 94 Vss 7.25701e-19
c142 89 Vss 9.96742e-19
c143 84 Vss 0.00258358f
c144 79 Vss 0.00309974f
c145 70 Vss 0.00527641f
c146 66 Vss 0.00738563f
c147 56 Vss 1.02723e-19
c148 54 Vss 0.0347733f
c149 53 Vss 0.0999357f
c150 42 Vss 0.035088f
c151 41 Vss 0.0994129f
c152 32 Vss 9.8832e-20
c153 30 Vss 0.0348822f
c154 29 Vss 0.10032f
c155 9 Vss 0.270154f
c156 7 Vss 0.269158f
c157 6 Vss 0.00143442f
c158 1 Vss 0.232685f
r159 149 161 0.494161
r160 149 151 6.54354
r161 145 161 0.128424
r162 144 160 0.494161
r163 143 155 0.652036
r164 143 144 7.46046
r165 139 160 0.128424
r166 137 161 0.494161
r167 137 138 15.8795
r168 133 159 0.0828784
r169 131 160 0.494161
r170 131 132 13.0037
r171 130 138 0.652036
r172 129 159 0.551426
r173 129 130 12.5036
r174 128 159 0.551426
r175 127 132 0.652036
r176 127 128 7.66886
r177 102 151 1.50043
r178 99 102 5.835
r179 94 119 1.16709
r180 94 155 2.16729
r181 89 114 1.16709
r182 89 145 2.16729
r183 84 139 5.2515
r184 79 105 1.16709
r185 79 133 4.33978
r186 70 99 1.16709
r187 66 84 1.16709
r188 56 119 0.0476429
r189 54 56 1.45875
r190 53 57 0.652036
r191 53 56 1.45875
r192 49 54 0.652036
r193 44 114 0.0476429
r194 42 44 1.45875
r195 41 45 0.652036
r196 41 44 1.45875
r197 37 42 0.652036
r198 32 105 0.238214
r199 30 32 1.45875
r200 29 33 0.652036
r201 29 32 1.45875
r202 25 30 0.652036
r203 12 70 0.185659
r204 9 57 3.8511
r205 9 49 3.8511
r206 7 45 3.8511
r207 7 37 3.8511
r208 6 66 0.185659
r209 4 66 0.185659
r210 1 33 3.1509
r211 1 25 3.1509
.ends

.subckt PM_G5_XNOR3_N2_CI 2 4 6 8 23 26 31 34 39 44 79 80 85 91 Vss
c48 91 Vss 2.53341e-19
c49 85 Vss 0.00608182f
c50 80 Vss 3.61784e-19
c51 79 Vss 0.00606729f
c52 44 Vss 0.00187346f
c53 39 Vss 0.00150573f
c54 34 Vss 0.00581447f
c55 31 Vss 0.00501461f
c56 26 Vss 0.00386883f
c57 23 Vss 0.00546807f
c58 4 Vss 0.00143442f
r59 86 91 0.441572
r60 85 87 0.655813
r61 85 86 9.04425
r62 81 91 0.174814
r63 79 91 0.441572
r64 79 80 19.1096
r65 75 80 0.655813
r66 44 87 2.41736
r67 39 81 2.41736
r68 34 75 13.4205
r69 31 44 1.16709
r70 26 39 1.16709
r71 23 34 1.16709
r72 8 31 0.185659
r73 6 26 0.185659
r74 4 23 0.185659
r75 2 23 0.185659
.ends

.subckt PM_G5_XNOR3_N2_A 2 4 5 7 20 44 45 49 55 58 60 61 66 69 70 73 78 Vss
c79 78 Vss 0.00548899f
c80 73 Vss 0.00489228f
c81 70 Vss 0.00566456f
c82 69 Vss 4.97253e-19
c83 61 Vss 5.64597e-19
c84 60 Vss 6.06847e-19
c85 58 Vss 0.00443885f
c86 55 Vss 0.00696223f
c87 49 Vss 0.135055f
c88 45 Vss 0.127825f
c89 44 Vss 9.8832e-20
c90 20 Vss 0.21515f
c91 17 Vss 0.129208f
c92 15 Vss 0.0247918f
c93 5 Vss 1.22081f
c94 4 Vss 0.139574f
r95 78 81 0.05
r96 69 81 1.16709
r97 69 70 0.531835
r98 64 73 1.16709
r99 64 66 0.125036
r100 61 64 0.833571
r101 60 70 10.4613
r102 57 60 0.652036
r103 57 58 8.66914
r104 56 61 0.0685365
r105 55 58 0.652036
r106 55 56 10.2113
r107 47 49 4.53833
r108 44 78 0.0238214
r109 44 45 2.26917
r110 41 44 2.26917
r111 34 49 0.00605528
r112 33 45 0.00605528
r113 28 47 0.00605528
r114 27 41 0.00605528
r115 23 73 0.0952857
r116 21 23 0.326018
r117 21 23 0.1167
r118 20 24 0.652036
r119 20 23 6.7686
r120 17 23 0.3335
r121 15 23 0.326018
r122 15 17 0.2334
r123 7 34 3.8511
r124 7 28 3.8511
r125 5 7 15.4044
r126 5 33 3.8511
r127 5 7 15.4044
r128 5 27 3.8511
r129 4 24 3.8511
r130 2 17 3.6177
.ends

.subckt PM_G5_XNOR3_N2_BI 2 4 6 8 16 23 29 32 37 42 51 56 64 65 71 77 82 83 Vss
c69 83 Vss 1.50773e-19
c70 82 Vss 0.00211439f
c71 77 Vss 0.00104035f
c72 71 Vss 3.29809e-19
c73 65 Vss 2.46443e-19
c74 64 Vss 0.00335376f
c75 56 Vss 0.00250661f
c76 51 Vss 0.00216609f
c77 42 Vss 0.00132272f
c78 37 Vss 9.45807e-19
c79 32 Vss 0.00229686f
c80 29 Vss 0.00450667f
c81 23 Vss 1.05854e-19
c82 16 Vss 0.111942f
c83 8 Vss 0.111942f
c84 4 Vss 0.00143442f
r85 81 83 0.65409
r86 81 82 3.42052
r87 77 82 0.652979
r88 64 71 0.0685365
r89 64 65 13.2121
r90 60 65 0.652036
r91 42 56 1.16709
r92 42 83 2.00578
r93 37 51 1.16709
r94 37 77 2.03284
r95 37 71 2.08393
r96 32 60 5.2515
r97 29 32 1.16709
r98 23 56 0.50025
r99 16 51 0.50025
r100 8 23 3.09255
r101 6 16 3.09255
r102 4 29 0.185659
r103 2 29 0.185659
.ends

.subckt PM_G5_XNOR3_N2_AI 2 4 5 7 31 37 43 50 55 64 72 Vss
c47 72 Vss 2.58509e-19
c48 64 Vss 0.005486f
c49 55 Vss 0.0041561f
c50 50 Vss 8.67602e-19
c51 43 Vss 0.00448756f
c52 37 Vss 0.127877f
c53 31 Vss 0.131783f
c54 5 Vss 1.2083f
c55 4 Vss 0.00143442f
r56 68 72 0.655813
r57 55 64 1.16709
r58 55 72 12.0347
r59 50 68 2.41736
r60 43 50 1.16709
r61 36 64 0.0238214
r62 36 37 2.334
r63 33 36 2.20433
r64 29 31 4.53833
r65 24 37 0.00605528
r66 23 31 0.00605528
r67 18 33 0.00605528
r68 17 29 0.00605528
r69 7 24 3.8511
r70 7 18 3.8511
r71 5 7 15.4044
r72 5 23 3.8511
r73 5 7 15.4044
r74 5 17 3.8511
r75 4 43 0.185659
r76 2 43 0.185659
.ends

.subckt PM_G5_XNOR3_N2_B 2 4 6 8 16 17 24 28 31 42 45 50 55 60 65 69 74 75 82
+ Vss
c65 82 Vss 3.53127e-19
c66 75 Vss 3.16204e-19
c67 74 Vss 7.66068e-19
c68 69 Vss 0.00368257f
c69 65 Vss 0.00255458f
c70 60 Vss 0.0023582f
c71 55 Vss 0.00157585f
c72 50 Vss 0.00115924f
c73 45 Vss 7.04295e-20
c74 42 Vss 5.36415e-19
c75 31 Vss 0.111942f
c76 24 Vss 1.02723e-19
c77 20 Vss 0.0247918f
c78 17 Vss 0.0338452f
c79 16 Vss 0.183686f
c80 6 Vss 0.112114f
c81 4 Vss 0.122719f
c82 2 Vss 0.13381f
r83 74 75 0.65409
r84 73 74 3.38028
r85 69 73 0.65409
r86 50 65 1.16709
r87 50 75 2.00578
r88 45 60 1.16709
r89 45 69 1.96931
r90 45 82 9.55481
r91 38 55 1.16709
r92 38 82 0.4602
r93 38 42 0.145875
r94 36 55 0.309679
r95 31 65 0.50025
r96 28 60 0.50025
r97 24 55 0.214393
r98 20 36 0.326018
r99 20 24 0.75855
r100 17 36 6.7686
r101 16 36 0.326018
r102 16 36 0.1167
r103 13 17 0.652036
r104 8 31 3.09255
r105 6 28 3.09255
r106 4 24 3.09255
r107 2 13 3.8511
.ends

.subckt PM_G5_XNOR3_N2_Z 2 4 6 8 23 27 30 33 Vss
c29 30 Vss 0.00359454f
c30 27 Vss 0.00857889f
c31 23 Vss 0.0074536f
c32 8 Vss 0.00143442f
c33 6 Vss 0.00143442f
r34 33 35 5.50157
r35 30 33 5.50157
r36 27 35 1.16709
r37 23 30 1.16709
r38 8 27 0.185659
r39 6 23 0.185659
r40 4 27 0.185659
r41 2 23 0.185659
.ends

.subckt G5_XNOR3_N2  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI13.X0 N_CI_XI13.X0_D N_VSS_XI13.X0_PGD N_C_XI13.X0_CG N_VSS_XI13.X0_PGD
+ N_VDD_XI13.X0_S TIGFET_HPNW8
XI16.X0 N_CI_XI16.X0_D N_VDD_XI16.X0_PGD N_C_XI16.X0_CG N_VDD_XI16.X0_PGD
+ N_VSS_XI16.X0_S TIGFET_HPNW8
XI15.X0 N_BI_XI15.X0_D N_VDD_XI15.X0_PGD N_B_XI15.X0_CG N_VDD_XI15.X0_PGD
+ N_VSS_XI15.X0_S TIGFET_HPNW8
XI11.X0 N_AI_XI11.X0_D N_VSS_XI11.X0_PGD N_A_XI11.X0_CG N_VSS_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW8
XI12.X0 N_BI_XI12.X0_D N_VSS_XI12.X0_PGD N_B_XI12.X0_CG N_VSS_XI12.X0_PGD
+ N_VDD_XI12.X0_S TIGFET_HPNW8
XI14.X0 N_AI_XI14.X0_D N_VDD_XI14.X0_PGD N_A_XI14.X0_CG N_VDD_XI14.X0_PGD
+ N_VSS_XI14.X0_S TIGFET_HPNW8
XI19.X0 N_Z_XI19.X0_D N_AI_XI19.X0_PGD N_B_XI19.X0_CG N_AI_XI19.X0_PGD
+ N_C_XI19.X0_S TIGFET_HPNW8
XI17.X0 N_Z_XI17.X0_D N_AI_XI17.X0_PGD N_BI_XI17.X0_CG N_AI_XI17.X0_PGD
+ N_CI_XI17.X0_S TIGFET_HPNW8
XI20.X0 N_Z_XI20.X0_D N_A_XI20.X0_PGD N_BI_XI20.X0_CG N_A_XI20.X0_PGD
+ N_C_XI20.X0_S TIGFET_HPNW8
XI18.X0 N_Z_XI18.X0_D N_A_XI18.X0_PGD N_B_XI18.X0_CG N_A_XI18.X0_PGD
+ N_CI_XI18.X0_S TIGFET_HPNW8
*
x_PM_G5_XNOR3_N2_VDD N_VDD_XI13.X0_S N_VDD_XI16.X0_PGD N_VDD_XI15.X0_PGD
+ N_VDD_XI11.X0_S N_VDD_XI12.X0_S N_VDD_XI14.X0_PGD N_VDD_c_115_p N_VDD_c_20_p
+ N_VDD_c_25_p N_VDD_c_3_p N_VDD_c_95_p N_VDD_c_106_p N_VDD_c_21_p N_VDD_c_77_p
+ N_VDD_c_107_p N_VDD_c_5_p N_VDD_c_6_p N_VDD_c_13_p N_VDD_c_4_p N_VDD_c_65_p
+ N_VDD_c_30_p N_VDD_c_66_p N_VDD_c_31_p N_VDD_c_17_p N_VDD_c_67_p N_VDD_c_22_p
+ N_VDD_c_10_p N_VDD_c_26_p N_VDD_c_38_p N_VDD_c_11_p N_VDD_c_61_p VDD
+ N_VDD_c_69_p N_VDD_c_73_p N_VDD_c_32_p N_VDD_c_43_p N_VDD_c_39_p Vss
+ PM_G5_XNOR3_N2_VDD
x_PM_G5_XNOR3_N2_C N_C_XI13.X0_CG N_C_XI16.X0_CG N_C_XI19.X0_S N_C_XI20.X0_S
+ N_C_c_118_n N_C_c_129_p N_C_c_121_n C N_C_c_122_n N_C_c_147_p N_C_c_144_p
+ N_C_c_124_n N_C_c_165_p N_C_c_126_n N_C_c_149_p N_C_c_154_p Vss
+ PM_G5_XNOR3_N2_C
x_PM_G5_XNOR3_N2_VSS N_VSS_XI13.X0_PGD N_VSS_XI16.X0_S N_VSS_XI15.X0_S
+ N_VSS_XI11.X0_PGD N_VSS_XI12.X0_PGD N_VSS_XI14.X0_S N_VSS_c_176_n
+ N_VSS_c_234_n N_VSS_c_177_n N_VSS_c_179_n N_VSS_c_180_n N_VSS_c_181_n
+ N_VSS_c_288_p N_VSS_c_183_n N_VSS_c_249_p N_VSS_c_184_n N_VSS_c_189_n
+ N_VSS_c_192_n N_VSS_c_196_n N_VSS_c_200_n N_VSS_c_203_n N_VSS_c_204_n
+ N_VSS_c_207_n N_VSS_c_211_n N_VSS_c_215_n N_VSS_c_218_n N_VSS_c_220_n
+ N_VSS_c_221_n N_VSS_c_222_n N_VSS_c_226_n N_VSS_c_227_n VSS N_VSS_c_230_n
+ N_VSS_c_231_n N_VSS_c_232_n Vss PM_G5_XNOR3_N2_VSS
x_PM_G5_XNOR3_N2_CI N_CI_XI13.X0_D N_CI_XI16.X0_D N_CI_XI17.X0_S N_CI_XI18.X0_S
+ N_CI_c_294_n N_CI_c_306_n N_CI_c_336_p N_CI_c_295_n N_CI_c_314_n N_CI_c_303_n
+ N_CI_c_299_n N_CI_c_319_n N_CI_c_322_p N_CI_c_331_p Vss PM_G5_XNOR3_N2_CI
x_PM_G5_XNOR3_N2_A N_A_XI11.X0_CG N_A_XI14.X0_CG N_A_XI20.X0_PGD N_A_XI18.X0_PGD
+ N_A_c_342_n N_A_c_376_p N_A_c_392_p N_A_c_394_p N_A_c_343_n N_A_c_349_n
+ N_A_c_350_n N_A_c_351_n A N_A_c_360_n N_A_c_361_n N_A_c_353_n N_A_c_382_p Vss
+ PM_G5_XNOR3_N2_A
x_PM_G5_XNOR3_N2_BI N_BI_XI15.X0_D N_BI_XI12.X0_D N_BI_XI17.X0_CG
+ N_BI_XI20.X0_CG N_BI_c_456_p N_BI_c_443_n N_BI_c_421_n N_BI_c_423_n
+ N_BI_c_459_p N_BI_c_438_n N_BI_c_457_p N_BI_c_450_n N_BI_c_427_n N_BI_c_454_n
+ N_BI_c_455_n N_BI_c_430_n N_BI_c_482_p N_BI_c_431_n Vss PM_G5_XNOR3_N2_BI
x_PM_G5_XNOR3_N2_AI N_AI_XI11.X0_D N_AI_XI14.X0_D N_AI_XI19.X0_PGD
+ N_AI_XI17.X0_PGD N_AI_c_499_n N_AI_c_491_n N_AI_c_492_n N_AI_c_494_n
+ N_AI_c_497_n N_AI_c_506_n N_AI_c_507_n Vss PM_G5_XNOR3_N2_AI
x_PM_G5_XNOR3_N2_B N_B_XI15.X0_CG N_B_XI12.X0_CG N_B_XI19.X0_CG N_B_XI18.X0_CG
+ N_B_c_538_n N_B_c_539_n N_B_c_545_n N_B_c_558_n N_B_c_559_n B N_B_c_562_n
+ N_B_c_551_n N_B_c_548_n N_B_c_567_n N_B_c_568_n N_B_c_540_n N_B_c_588_n
+ N_B_c_552_n N_B_c_550_n Vss PM_G5_XNOR3_N2_B
x_PM_G5_XNOR3_N2_Z N_Z_XI19.X0_D N_Z_XI17.X0_D N_Z_XI20.X0_D N_Z_XI18.X0_D
+ N_Z_c_602_n N_Z_c_608_n N_Z_c_606_n Z Vss PM_G5_XNOR3_N2_Z
cc_1 N_VDD_XI15.X0_PGD N_C_XI16.X0_CG 0.00111638f
cc_2 N_VDD_XI16.X0_PGD N_C_c_118_n 4.18107e-19
cc_3 N_VDD_c_3_p N_C_c_118_n 0.00111638f
cc_4 N_VDD_c_4_p N_C_c_118_n 0.00134502f
cc_5 N_VDD_c_5_p N_C_c_121_n 3.43419e-19
cc_6 N_VDD_c_6_p N_C_c_122_n 4.34606e-19
cc_7 N_VDD_c_4_p N_C_c_122_n 0.00156986f
cc_8 N_VDD_c_6_p N_C_c_124_n 4.60895e-19
cc_9 N_VDD_c_4_p N_C_c_124_n 2.85335e-19
cc_10 N_VDD_c_10_p N_C_c_126_n 4.68396e-19
cc_11 N_VDD_c_11_p N_C_c_126_n 7.76004e-19
cc_12 N_VDD_XI16.X0_PGD N_VSS_XI13.X0_PGD 0.00162006f
cc_13 N_VDD_c_13_p N_VSS_XI13.X0_PGD 2.10457e-19
cc_14 N_VDD_c_4_p N_VSS_XI13.X0_PGD 2.00345e-19
cc_15 N_VDD_XI15.X0_PGD N_VSS_XI11.X0_PGD 2.37403e-19
cc_16 N_VDD_XI14.X0_PGD N_VSS_XI11.X0_PGD 0.00200476f
cc_17 N_VDD_c_17_p N_VSS_XI11.X0_PGD 2.94729e-19
cc_18 N_VDD_XI15.X0_PGD N_VSS_XI12.X0_PGD 0.00200584f
cc_19 N_VDD_XI14.X0_PGD N_VSS_XI12.X0_PGD 2.24644e-19
cc_20 N_VDD_c_20_p N_VSS_c_176_n 0.00162006f
cc_21 N_VDD_c_21_p N_VSS_c_177_n 0.00200476f
cc_22 N_VDD_c_22_p N_VSS_c_177_n 2.84318e-19
cc_23 N_VDD_c_22_p N_VSS_c_179_n 3.9313e-19
cc_24 N_VDD_c_11_p N_VSS_c_180_n 2.35523e-19
cc_25 N_VDD_c_25_p N_VSS_c_181_n 0.00200584f
cc_26 N_VDD_c_26_p N_VSS_c_181_n 3.9313e-19
cc_27 N_VDD_c_4_p N_VSS_c_183_n 3.4118e-19
cc_28 N_VDD_c_13_p N_VSS_c_184_n 4.32468e-19
cc_29 N_VDD_c_4_p N_VSS_c_184_n 4.11891e-19
cc_30 N_VDD_c_30_p N_VSS_c_184_n 0.00126261f
cc_31 N_VDD_c_31_p N_VSS_c_184_n 3.98949e-19
cc_32 N_VDD_c_32_p N_VSS_c_184_n 3.48267e-19
cc_33 N_VDD_c_4_p N_VSS_c_189_n 3.98099e-19
cc_34 N_VDD_c_10_p N_VSS_c_189_n 7.41581e-19
cc_35 N_VDD_c_11_p N_VSS_c_189_n 5.12345e-19
cc_36 N_VDD_c_17_p N_VSS_c_192_n 6.9475e-19
cc_37 N_VDD_c_22_p N_VSS_c_192_n 0.00161703f
cc_38 N_VDD_c_38_p N_VSS_c_192_n 9.10421e-19
cc_39 N_VDD_c_39_p N_VSS_c_192_n 3.48267e-19
cc_40 N_VDD_c_10_p N_VSS_c_196_n 6.80981e-19
cc_41 N_VDD_c_26_p N_VSS_c_196_n 0.00161703f
cc_42 N_VDD_c_11_p N_VSS_c_196_n 0.00260511f
cc_43 N_VDD_c_43_p N_VSS_c_196_n 3.48267e-19
cc_44 N_VDD_XI14.X0_PGD N_VSS_c_200_n 2.99706e-19
cc_45 N_VDD_c_38_p N_VSS_c_200_n 0.00524008f
cc_46 N_VDD_c_39_p N_VSS_c_200_n 9.58524e-19
cc_47 N_VDD_c_22_p N_VSS_c_203_n 0.00398219f
cc_48 N_VDD_c_13_p N_VSS_c_204_n 4.41003e-19
cc_49 N_VDD_c_31_p N_VSS_c_204_n 3.89161e-19
cc_50 N_VDD_c_32_p N_VSS_c_204_n 6.39485e-19
cc_51 N_VDD_c_17_p N_VSS_c_207_n 3.48267e-19
cc_52 N_VDD_c_22_p N_VSS_c_207_n 2.26455e-19
cc_53 N_VDD_c_38_p N_VSS_c_207_n 3.99794e-19
cc_54 N_VDD_c_39_p N_VSS_c_207_n 6.489e-19
cc_55 N_VDD_c_10_p N_VSS_c_211_n 3.82294e-19
cc_56 N_VDD_c_26_p N_VSS_c_211_n 2.26455e-19
cc_57 N_VDD_c_11_p N_VSS_c_211_n 9.55109e-19
cc_58 N_VDD_c_43_p N_VSS_c_211_n 6.46219e-19
cc_59 N_VDD_c_6_p N_VSS_c_215_n 0.00346699f
cc_60 N_VDD_c_13_p N_VSS_c_215_n 0.0014056f
cc_61 N_VDD_c_61_p N_VSS_c_215_n 0.0010705f
cc_62 N_VDD_c_13_p N_VSS_c_218_n 0.00935412f
cc_63 N_VDD_c_31_p N_VSS_c_218_n 0.00107899f
cc_64 N_VDD_c_4_p N_VSS_c_220_n 0.00942626f
cc_65 N_VDD_c_65_p N_VSS_c_221_n 0.00107364f
cc_66 N_VDD_c_66_p N_VSS_c_222_n 0.00824191f
cc_67 N_VDD_c_67_p N_VSS_c_222_n 7.27535e-19
cc_68 N_VDD_c_22_p N_VSS_c_222_n 0.00364308f
cc_69 N_VDD_c_69_p N_VSS_c_222_n 0.00146091f
cc_70 N_VDD_c_13_p N_VSS_c_226_n 0.00107577f
cc_71 N_VDD_c_4_p N_VSS_c_227_n 0.00143205f
cc_72 N_VDD_c_26_p N_VSS_c_227_n 0.00595362f
cc_73 N_VDD_c_73_p N_VSS_c_227_n 0.00107225f
cc_74 N_VDD_c_13_p N_VSS_c_230_n 0.00112682f
cc_75 N_VDD_c_4_p N_VSS_c_231_n 0.00107375f
cc_76 N_VDD_c_22_p N_VSS_c_232_n 7.74609e-19
cc_77 N_VDD_c_77_p N_CI_c_294_n 3.43419e-19
cc_78 N_VDD_c_77_p N_CI_c_295_n 3.48267e-19
cc_79 N_VDD_c_4_p N_CI_c_295_n 4.34701e-19
cc_80 N_VDD_c_30_p N_CI_c_295_n 5.61123e-19
cc_81 N_VDD_c_31_p N_CI_c_295_n 0.00251349f
cc_82 N_VDD_c_17_p N_CI_c_299_n 9.69348e-19
cc_83 N_VDD_c_67_p N_CI_c_299_n 5.49852e-19
cc_84 N_VDD_XI14.X0_PGD N_A_c_342_n 3.94724e-19
cc_85 N_VDD_XI14.X0_PGD N_A_c_343_n 4.9801e-19
cc_86 N_VDD_c_5_p N_A_c_343_n 2.69869e-19
cc_87 N_VDD_c_22_p N_A_c_343_n 2.92916e-19
cc_88 N_VDD_c_38_p N_A_c_343_n 2.57998e-19
cc_89 N_VDD_c_11_p N_A_c_343_n 3.18391e-19
cc_90 N_VDD_c_39_p N_A_c_343_n 4.99558e-19
cc_91 N_VDD_c_5_p N_A_c_349_n 9.18655e-19
cc_92 N_VDD_c_11_p N_A_c_350_n 0.00561464f
cc_93 N_VDD_c_31_p N_A_c_351_n 0.00109781f
cc_94 N_VDD_c_10_p N_A_c_351_n 2.35756e-19
cc_95 N_VDD_c_95_p N_A_c_353_n 3.65048e-19
cc_96 N_VDD_c_31_p N_A_c_353_n 5.7233e-19
cc_97 N_VDD_c_43_p N_A_c_353_n 2.01103e-19
cc_98 N_VDD_c_5_p N_BI_c_421_n 3.43419e-19
cc_99 N_VDD_c_11_p N_BI_c_421_n 3.48267e-19
cc_100 N_VDD_c_5_p N_BI_c_423_n 3.48267e-19
cc_101 N_VDD_c_31_p N_BI_c_423_n 9.37844e-19
cc_102 N_VDD_c_26_p N_BI_c_423_n 4.34701e-19
cc_103 N_VDD_c_11_p N_BI_c_423_n 4.99861e-19
cc_104 N_VDD_c_26_p N_BI_c_427_n 2.93466e-19
cc_105 N_VDD_XI14.X0_PGD N_AI_XI19.X0_PGD 3.10667e-19
cc_106 N_VDD_c_106_p N_AI_c_491_n 3.10667e-19
cc_107 N_VDD_c_107_p N_AI_c_492_n 3.43419e-19
cc_108 N_VDD_c_67_p N_AI_c_492_n 3.73302e-19
cc_109 N_VDD_c_107_p N_AI_c_494_n 3.48267e-19
cc_110 N_VDD_c_67_p N_AI_c_494_n 5.23123e-19
cc_111 N_VDD_c_22_p N_AI_c_494_n 4.34701e-19
cc_112 N_VDD_c_38_p N_AI_c_497_n 0.00114561f
cc_113 N_VDD_XI16.X0_PGD N_B_XI15.X0_CG 8.43351e-19
cc_114 N_VDD_XI15.X0_PGD N_B_c_538_n 3.99339e-19
cc_115 N_VDD_c_115_p N_B_c_539_n 8.43351e-19
cc_116 N_VDD_c_11_p N_B_c_540_n 4.93279e-19
cc_117 N_C_c_118_n N_VSS_XI13.X0_PGD 4.18107e-19
cc_118 N_C_c_129_p N_VSS_c_234_n 9.69352e-19
cc_119 N_C_c_122_n N_VSS_c_184_n 7.02166e-19
cc_120 N_C_c_124_n N_VSS_c_184_n 3.26762e-19
cc_121 N_C_c_122_n N_VSS_c_189_n 2.08725e-19
cc_122 N_C_c_126_n N_VSS_c_189_n 0.00161414f
cc_123 N_C_c_126_n N_VSS_c_196_n 0.00142183f
cc_124 N_C_c_122_n N_VSS_c_204_n 3.26762e-19
cc_125 N_C_c_124_n N_VSS_c_204_n 2.75266e-19
cc_126 N_C_c_122_n N_VSS_c_215_n 4.20305e-19
cc_127 N_C_c_126_n N_VSS_c_215_n 2.33946e-19
cc_128 N_C_c_122_n N_VSS_c_220_n 0.00170504f
cc_129 N_C_c_126_n N_VSS_c_220_n 0.00306503f
cc_130 N_C_c_126_n N_VSS_c_227_n 0.00185247f
cc_131 N_C_c_118_n N_CI_c_294_n 6.55689e-19
cc_132 N_C_c_126_n N_CI_c_295_n 0.00101197f
cc_133 N_C_c_144_p N_CI_c_303_n 2.42706e-19
cc_134 N_C_c_126_n N_A_c_343_n 3.07864e-19
cc_135 N_C_c_121_n N_A_c_349_n 8.20481e-19
cc_136 N_C_c_147_p N_A_c_349_n 0.00174813f
cc_137 N_C_c_126_n N_A_c_350_n 3.74205e-19
cc_138 N_C_c_149_p N_A_c_360_n 3.98753e-19
cc_139 N_C_c_121_n N_A_c_361_n 8.20481e-19
cc_140 N_C_c_147_p N_A_c_361_n 0.00170439f
cc_141 N_C_c_126_n N_A_c_361_n 3.354e-19
cc_142 N_C_c_149_p N_A_c_361_n 0.00192636f
cc_143 N_C_c_154_p N_A_c_361_n 2.01694e-19
cc_144 N_C_c_126_n N_BI_c_423_n 4.79207e-19
cc_145 N_C_c_126_n N_BI_c_427_n 5.14704e-19
cc_146 N_C_c_149_p N_BI_c_430_n 5.49277e-19
cc_147 N_C_c_149_p N_BI_c_431_n 0.00181681f
cc_148 N_C_c_147_p N_B_c_540_n 0.00168209f
cc_149 N_C_c_126_n N_B_c_540_n 0.00270379f
cc_150 N_C_c_149_p N_B_c_540_n 0.0010597f
cc_151 N_C_c_121_n N_Z_c_602_n 3.43419e-19
cc_152 N_C_c_147_p N_Z_c_602_n 3.48267e-19
cc_153 N_C_c_144_p N_Z_c_602_n 3.48267e-19
cc_154 N_C_c_165_p N_Z_c_602_n 3.43419e-19
cc_155 N_C_c_147_p N_Z_c_606_n 6.10113e-19
cc_156 N_C_c_144_p N_Z_c_606_n 5.74072e-19
cc_157 N_VSS_c_183_n N_CI_c_294_n 3.43419e-19
cc_158 N_VSS_c_189_n N_CI_c_294_n 3.48267e-19
cc_159 N_VSS_c_249_p N_CI_c_306_n 3.43419e-19
cc_160 N_VSS_c_200_n N_CI_c_306_n 3.48267e-19
cc_161 N_VSS_c_183_n N_CI_c_295_n 3.48267e-19
cc_162 N_VSS_c_184_n N_CI_c_295_n 5.78167e-19
cc_163 N_VSS_c_189_n N_CI_c_295_n 0.00107566f
cc_164 N_VSS_c_215_n N_CI_c_295_n 3.18991e-19
cc_165 N_VSS_c_218_n N_CI_c_295_n 0.00247956f
cc_166 N_VSS_c_220_n N_CI_c_295_n 2.82247e-19
cc_167 N_VSS_c_249_p N_CI_c_314_n 3.48267e-19
cc_168 N_VSS_c_200_n N_CI_c_314_n 9.64594e-19
cc_169 N_VSS_c_192_n N_CI_c_299_n 0.00118348f
cc_170 N_VSS_c_203_n N_CI_c_299_n 0.0033401f
cc_171 N_VSS_c_222_n N_CI_c_299_n 2.16087e-19
cc_172 N_VSS_c_222_n N_CI_c_319_n 0.00291606f
cc_173 N_VSS_XI11.X0_PGD N_A_c_342_n 3.91527e-19
cc_174 N_VSS_c_249_p N_A_c_343_n 5.38503e-19
cc_175 N_VSS_c_200_n N_A_c_343_n 8.92829e-19
cc_176 N_VSS_c_203_n N_A_c_343_n 2.86582e-19
cc_177 N_VSS_c_192_n N_A_c_351_n 3.11664e-19
cc_178 N_VSS_c_207_n N_A_c_351_n 3.1261e-19
cc_179 N_VSS_c_192_n N_A_c_353_n 3.04912e-19
cc_180 N_VSS_c_207_n N_A_c_353_n 0.00110478f
cc_181 N_VSS_c_183_n N_BI_c_421_n 3.43419e-19
cc_182 N_VSS_c_189_n N_BI_c_421_n 3.48267e-19
cc_183 N_VSS_c_183_n N_BI_c_423_n 3.48267e-19
cc_184 N_VSS_c_189_n N_BI_c_423_n 0.00102079f
cc_185 N_VSS_c_227_n N_BI_c_423_n 2.89128e-19
cc_186 N_VSS_XI12.X0_PGD N_AI_XI19.X0_PGD 2.79882e-19
cc_187 N_VSS_c_180_n N_AI_c_499_n 2.79882e-19
cc_188 N_VSS_c_249_p N_AI_c_492_n 3.43419e-19
cc_189 N_VSS_c_200_n N_AI_c_492_n 3.48267e-19
cc_190 N_VSS_c_249_p N_AI_c_494_n 3.48267e-19
cc_191 N_VSS_c_200_n N_AI_c_494_n 0.001398f
cc_192 N_VSS_c_200_n N_AI_c_497_n 0.00172519f
cc_193 N_VSS_c_203_n N_AI_c_497_n 0.00643151f
cc_194 N_VSS_c_200_n N_AI_c_506_n 2.82216e-19
cc_195 N_VSS_c_192_n N_AI_c_507_n 0.00195338f
cc_196 N_VSS_c_203_n N_AI_c_507_n 0.00167155f
cc_197 N_VSS_XI12.X0_PGD N_B_c_538_n 3.96142e-19
cc_198 N_VSS_c_288_p N_B_c_545_n 0.00112923f
cc_199 N_VSS_c_196_n B 3.70276e-19
cc_200 N_VSS_c_211_n B 3.65807e-19
cc_201 N_VSS_c_196_n N_B_c_548_n 3.65807e-19
cc_202 N_VSS_c_211_n N_B_c_548_n 3.61194e-19
cc_203 N_VSS_c_196_n N_B_c_550_n 4.74612e-19
cc_204 N_CI_c_299_n N_A_c_343_n 4.46962e-19
cc_205 N_CI_c_295_n N_BI_c_423_n 0.00125164f
cc_206 N_CI_c_322_p N_BI_c_438_n 6.43262e-19
cc_207 N_CI_c_314_n N_BI_c_427_n 5.16242e-19
cc_208 N_CI_c_299_n N_BI_c_427_n 0.00141805f
cc_209 N_CI_c_322_p N_BI_c_430_n 0.00184196f
cc_210 N_CI_c_295_n N_AI_c_494_n 5.9142e-19
cc_211 N_CI_c_314_n N_AI_c_494_n 5.87215e-19
cc_212 N_CI_c_314_n N_AI_c_497_n 0.00175375f
cc_213 N_CI_c_299_n N_AI_c_497_n 0.0058239f
cc_214 N_CI_c_322_p N_AI_c_497_n 0.00302067f
cc_215 N_CI_c_331_p N_AI_c_497_n 9.17939e-19
cc_216 N_CI_c_299_n N_AI_c_507_n 6.9086e-19
cc_217 N_CI_c_322_p N_B_c_551_n 8.97242e-19
cc_218 N_CI_c_322_p N_B_c_552_n 2.22052e-19
cc_219 N_CI_c_306_n N_Z_c_608_n 3.43419e-19
cc_220 N_CI_c_336_p N_Z_c_608_n 3.43419e-19
cc_221 N_CI_c_314_n N_Z_c_608_n 3.48267e-19
cc_222 N_CI_c_303_n N_Z_c_608_n 3.48267e-19
cc_223 N_CI_c_336_p N_Z_c_606_n 3.48267e-19
cc_224 N_CI_c_314_n N_Z_c_606_n 6.09821e-19
cc_225 N_CI_c_303_n N_Z_c_606_n 5.71987e-19
cc_226 N_A_XI20.X0_PGD N_BI_XI20.X0_CG 9.65637e-19
cc_227 N_A_c_376_p N_BI_c_443_n 9.50932e-19
cc_228 N_A_c_343_n N_BI_c_421_n 2.69869e-19
cc_229 N_A_c_343_n N_BI_c_423_n 2.84781e-19
cc_230 N_A_c_349_n N_BI_c_423_n 7.93978e-19
cc_231 N_A_c_360_n N_BI_c_438_n 5.59762e-19
cc_232 N_A_c_361_n N_BI_c_438_n 2.11253e-19
cc_233 N_A_c_382_p N_BI_c_438_n 3.26762e-19
cc_234 N_A_XI20.X0_PGD N_BI_c_450_n 0.00133285f
cc_235 N_A_c_382_p N_BI_c_450_n 2.75266e-19
cc_236 N_A_c_343_n N_BI_c_427_n 0.0032866f
cc_237 N_A_c_349_n N_BI_c_427_n 0.00143358f
cc_238 N_A_c_343_n N_BI_c_454_n 6.46327e-19
cc_239 N_A_c_343_n N_BI_c_455_n 2.29103e-19
cc_240 N_A_XI20.X0_PGD N_AI_XI19.X0_PGD 0.0174153f
cc_241 N_A_c_349_n N_AI_XI19.X0_PGD 9.9436e-19
cc_242 N_A_c_361_n N_AI_XI19.X0_PGD 0.00100436f
cc_243 N_A_c_392_p N_AI_c_499_n 0.00199603f
cc_244 N_A_c_361_n N_AI_c_499_n 0.001261f
cc_245 N_A_c_394_p N_AI_c_491_n 0.00201004f
cc_246 N_A_c_342_n N_AI_c_492_n 6.8653e-19
cc_247 N_A_c_343_n N_AI_c_494_n 8.04759e-19
cc_248 N_A_c_343_n N_AI_c_497_n 0.00144224f
cc_249 N_A_c_342_n N_B_c_538_n 0.00359928f
cc_250 N_A_c_343_n N_B_c_538_n 3.71868e-19
cc_251 N_A_c_351_n N_B_c_539_n 3.71868e-19
cc_252 N_A_c_353_n N_B_c_539_n 5.91713e-19
cc_253 N_A_c_343_n N_B_c_545_n 3.88197e-19
cc_254 N_A_c_361_n N_B_c_558_n 2.74063e-19
cc_255 N_A_XI20.X0_PGD N_B_c_559_n 9.65637e-19
cc_256 N_A_c_343_n B 7.21228e-19
cc_257 N_A_c_349_n B 4.92712e-19
cc_258 N_A_c_349_n N_B_c_562_n 3.80412e-19
cc_259 N_A_c_361_n N_B_c_562_n 3.68965e-19
cc_260 N_A_c_361_n N_B_c_551_n 4.34114e-19
cc_261 N_A_c_342_n N_B_c_548_n 6.98561e-19
cc_262 N_A_c_349_n N_B_c_548_n 6.04163e-19
cc_263 N_A_c_349_n N_B_c_567_n 3.37713e-19
cc_264 N_A_XI20.X0_PGD N_B_c_568_n 0.00133285f
cc_265 N_A_c_343_n N_B_c_540_n 0.00124487f
cc_266 N_A_c_349_n N_B_c_540_n 0.00208788f
cc_267 N_A_c_361_n N_B_c_540_n 0.00263274f
cc_268 N_A_c_361_n N_Z_c_602_n 0.00109616f
cc_269 N_A_XI20.X0_PGD N_Z_c_606_n 7.88059e-19
cc_270 N_A_c_349_n N_Z_c_606_n 0.00136894f
cc_271 N_A_c_361_n N_Z_c_606_n 0.00142189f
cc_272 N_BI_c_456_p N_AI_XI19.X0_PGD 9.65637e-19
cc_273 N_BI_c_457_p N_AI_XI19.X0_PGD 0.00133285f
cc_274 N_BI_c_454_n N_AI_c_494_n 5.87796e-19
cc_275 N_BI_c_459_p N_AI_c_497_n 3.22026e-19
cc_276 N_BI_c_457_p N_AI_c_497_n 3.2351e-19
cc_277 N_BI_c_427_n N_AI_c_497_n 0.00274992f
cc_278 N_BI_c_455_n N_AI_c_497_n 2.49817e-19
cc_279 N_BI_c_459_p N_AI_c_506_n 3.26631e-19
cc_280 N_BI_c_457_p N_AI_c_506_n 0.00116273f
cc_281 N_BI_c_421_n N_B_c_538_n 6.8653e-19
cc_282 N_BI_c_423_n B 4.49325e-19
cc_283 N_BI_c_459_p N_B_c_562_n 6.00485e-19
cc_284 N_BI_c_457_p N_B_c_562_n 4.7755e-19
cc_285 N_BI_c_455_n N_B_c_562_n 3.12886e-19
cc_286 N_BI_c_438_n N_B_c_551_n 0.00178472f
cc_287 N_BI_c_459_p N_B_c_567_n 4.95293e-19
cc_288 N_BI_c_457_p N_B_c_567_n 0.00384234f
cc_289 N_BI_c_450_n N_B_c_567_n 6.17967e-19
cc_290 N_BI_c_438_n N_B_c_568_n 4.56568e-19
cc_291 N_BI_c_457_p N_B_c_568_n 7.16621e-19
cc_292 N_BI_c_450_n N_B_c_568_n 0.00243716f
cc_293 N_BI_c_438_n N_B_c_540_n 0.00166188f
cc_294 N_BI_c_455_n N_B_c_540_n 0.0081489f
cc_295 N_BI_c_430_n N_B_c_540_n 7.19198e-19
cc_296 N_BI_c_431_n N_B_c_540_n 8.87908e-19
cc_297 N_BI_c_455_n N_B_c_588_n 0.00345251f
cc_298 N_BI_c_482_p N_B_c_588_n 0.00190039f
cc_299 N_BI_c_430_n N_B_c_552_n 8.29167e-19
cc_300 N_BI_c_423_n N_B_c_550_n 0.00221197f
cc_301 N_BI_c_427_n N_B_c_550_n 0.0081489f
cc_302 N_BI_c_459_p N_Z_c_606_n 0.00181417f
cc_303 N_BI_c_438_n N_Z_c_606_n 0.00138952f
cc_304 N_BI_c_450_n N_Z_c_606_n 8.66889e-19
cc_305 N_BI_c_455_n N_Z_c_606_n 4.80971e-19
cc_306 N_AI_XI19.X0_PGD N_B_XI19.X0_CG 9.47088e-19
cc_307 N_AI_XI19.X0_PGD N_B_c_567_n 0.00133285f
cc_308 N_AI_XI19.X0_PGD N_Z_c_606_n 4.24145e-19
cc_309 N_B_c_562_n N_Z_c_606_n 0.00138952f
cc_310 N_B_c_551_n N_Z_c_606_n 0.00138952f
cc_311 N_B_c_567_n N_Z_c_606_n 8.66889e-19
cc_312 N_B_c_568_n N_Z_c_606_n 8.66889e-19
cc_313 N_B_c_540_n N_Z_c_606_n 0.0010571f
cc_314 N_B_c_588_n N_Z_c_606_n 0.00213616f
cc_315 N_B_c_552_n N_Z_c_606_n 0.00102447f
*
.ends
*
*
.subckt XNOR3_HPNW8 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XNOR3_N2
.ends
*
* File: G4_XOR2_N2.pex.netlist
* Created: Sun Apr 10 19:56:43 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XOR2_N2_VSS 2 5 9 12 14 16 32 33 42 43 45 54 59 63 66 71 76 81 86
+ 95 100 113 115 116 117 122 123 128 138 140 145 146 147 150
c98 148 0 6.15603e-19
c99 147 0 3.75522e-19
c100 146 0 4.28045e-19
c101 145 0 0.00386476f
c102 140 0 0.0021378f
c103 138 0 0.00844222f
c104 128 0 0.00339884f
c105 123 0 8.42592e-19
c106 122 0 0.00171246f
c107 117 0 8.20625e-19
c108 116 0 0.00418359f
c109 115 0 0.00524404f
c110 113 0 0.00159018f
c111 100 0 0.00404792f
c112 95 0 0.00404489f
c113 86 0 1.66825e-19
c114 81 0 0.00174451f
c115 76 0 6.28678e-19
c116 71 0 9.88359e-19
c117 66 0 0.00180488f
c118 63 0 0.00552459f
c119 59 0 0.00736499f
c120 54 0 0.00542864f
c121 45 0 1.03318e-19
c122 43 0 0.0342891f
c123 42 0 0.100068f
c124 33 0 0.0350852f
c125 32 0 0.0990727f
c126 14 0 0.00143442f
c127 9 0 0.269235f
c128 5 0 0.268907f
r129 145 150 0.326018
r130 144 145 4.58464
r131 140 144 0.655813
r132 139 148 0.494161
r133 138 150 0.326018
r134 138 139 13.0037
r135 134 148 0.128424
r136 129 147 0.494161
r137 128 148 0.494161
r138 128 129 7.46046
r139 124 147 0.128424
r140 122 147 0.494161
r141 122 123 4.37625
r142 118 146 0.0828784
r143 116 130 0.652036
r144 116 117 10.1279
r145 115 123 0.652036
r146 114 146 0.551426
r147 114 115 14.4208
r148 113 146 0.551426
r149 112 117 0.652036
r150 112 113 4.58464
r151 86 140 1.82344
r152 81 134 5.2515
r153 76 100 1.16709
r154 76 130 2.16729
r155 71 95 1.16709
r156 71 124 2.16729
r157 66 118 1.82344
r158 63 86 1.16709
r159 59 81 1.16709
r160 54 66 1.16709
r161 45 100 0.0476429
r162 43 45 1.45875
r163 42 46 0.652036
r164 42 45 1.45875
r165 39 43 0.652036
r166 35 95 0.0476429
r167 33 35 1.45875
r168 32 36 0.652036
r169 32 35 1.45875
r170 29 33 0.652036
r171 16 63 0.185659
r172 14 59 0.185659
r173 12 59 0.185659
r174 9 46 3.8511
r175 9 39 3.8511
r176 5 36 3.8511
r177 5 29 3.8511
r178 2 54 0.185659
.ends

.subckt PM_G4_XOR2_N2_VDD 3 6 8 11 14 16 32 42 43 54 59 63 66 68 69 70 73 75 76
+ 79 81 85 89 91 93 98 99 100 103 109 114
c99 114 0 0.00454282f
c100 109 0 0.00472544f
c101 101 0 8.79456e-19
c102 100 0 2.39889e-19
c103 99 0 4.52364e-19
c104 98 0 0.00483655f
c105 93 0 0.00147365f
c106 91 0 0.0130047f
c107 89 0 0.00227129f
c108 85 0 8.26969e-19
c109 81 0 0.00455615f
c110 79 0 0.00100252f
c111 76 0 8.63853e-19
c112 75 0 0.0057282f
c113 73 0 0.0019575f
c114 70 0 8.67926e-19
c115 69 0 0.00221146f
c116 68 0 0.00205498f
c117 66 0 0.00803904f
c118 63 0 0.00389115f
c119 59 0 0.00739215f
c120 54 0 0.00398638f
c121 43 0 0.0351228f
c122 42 0 0.100954f
c123 35 0 2.09107e-19
c124 33 0 0.035919f
c125 32 0 0.100953f
c126 14 0 0.00143442f
c127 11 0 0.269396f
c128 3 0 0.270542f
r129 98 103 0.349767
r130 97 98 4.58464
r131 93 103 0.306046
r132 93 95 1.82344
r133 92 101 0.494161
r134 91 97 0.652036
r135 91 92 13.0037
r136 87 101 0.128424
r137 87 89 5.2515
r138 85 114 1.16709
r139 83 85 2.16729
r140 82 100 0.494161
r141 81 101 0.494161
r142 81 82 7.46046
r143 79 109 1.16709
r144 77 100 0.128424
r145 77 79 2.16729
r146 75 83 0.652036
r147 75 76 10.1279
r148 71 99 0.0828784
r149 71 73 1.82344
r150 69 100 0.494161
r151 69 70 4.37625
r152 68 76 0.652036
r153 67 99 0.551426
r154 67 68 4.58464
r155 66 99 0.551426
r156 65 70 0.652036
r157 65 66 14.4208
r158 63 95 1.16709
r159 59 89 1.16709
r160 54 73 1.02121
r161 45 114 0.0476429
r162 43 45 1.45875
r163 42 46 0.652036
r164 42 45 1.45875
r165 39 43 0.652036
r166 35 109 0.0476429
r167 33 35 1.45875
r168 32 36 0.652036
r169 32 35 1.45875
r170 29 33 0.652036
r171 16 63 0.185659
r172 14 59 0.185659
r173 11 46 3.8511
r174 11 39 3.8511
r175 8 59 0.185659
r176 6 54 0.185659
r177 3 36 3.8511
r178 3 29 3.8511
.ends

.subckt PM_G4_XOR2_N2_A 2 4 7 10 21 24 28 39 48 51 54 57 62 67 72 77 85
c58 85 0 8.29046e-19
c59 77 0 0.00201173f
c60 72 0 0.00648506f
c61 67 0 0.00351476f
c62 62 0 0.00246599f
c63 57 0 0.00406665f
c64 54 0 7.62653e-19
c65 48 0 0.128037f
c66 43 0 0.0296312f
c67 39 0 2.38608e-19
c68 28 0 0.152668f
c69 24 0 9.84889e-20
c70 21 0 0.169628f
c71 18 0 0.126125f
c72 16 0 0.0247918f
c73 10 0 0.1218f
c74 7 0 0.324846f
c75 4 0 0.138512f
r76 81 85 0.653045
r77 62 77 1.16709
r78 62 85 4.9014
r79 57 72 1.16709
r80 57 81 9.00257
r81 54 67 1.16709
r82 51 54 0.0364688
r83 47 72 0.0238214
r84 47 48 2.334
r85 44 47 2.20433
r86 39 77 0.50025
r87 33 48 0.00605528
r88 31 44 0.00605528
r89 29 43 0.494161
r90 28 30 0.652036
r91 28 29 4.84305
r92 25 43 0.128424
r93 24 67 0.0476429
r94 22 24 0.326018
r95 22 24 0.1167
r96 21 43 0.494161
r97 21 24 6.7686
r98 18 67 0.357321
r99 16 24 0.326018
r100 16 18 0.40845
r101 10 39 3.3843
r102 7 33 3.8511
r103 7 31 3.8511
r104 7 30 3.8511
r105 4 25 3.8511
r106 2 18 3.44265
.ends

.subckt PM_G4_XOR2_N2_NET1 2 4 7 10 30 31 35 41 44 49 58 76
c37 76 0 3.4517e-19
c38 58 0 0.00413905f
c39 49 0 0.00667491f
c40 44 0 0.00198364f
c41 41 0 0.00539823f
c42 35 0 0.103124f
c43 31 0 0.125482f
c44 30 0 9.62407e-20
c45 10 0 0.214624f
c46 7 0 0.384182f
c47 4 0 0.00143442f
r48 72 76 0.655813
r49 49 58 1.16709
r50 49 76 12.1076
r51 44 72 2.41736
r52 41 44 1.16709
r53 33 35 1.70187
r54 30 58 0.0238214
r55 30 31 2.20433
r56 27 30 2.334
r57 25 35 0.17282
r58 24 31 0.00605528
r59 21 33 0.17282
r60 18 27 0.00605528
r61 10 21 6.36015
r62 7 25 6.01005
r63 7 24 3.8511
r64 7 18 3.8511
r65 4 41 0.185659
r66 2 41 0.185659
.ends

.subckt PM_G4_XOR2_N2_NET2 2 4 6 9 21 22 33 39 42 47 56 74
c44 74 0 3.04338e-19
c45 56 0 0.00509819f
c46 47 0 0.00799947f
c47 42 0 0.00221316f
c48 39 0 0.00534974f
c49 33 0 0.129063f
c50 22 0 0.0345383f
c51 21 0 0.17396f
c52 9 0 0.466016f
c53 6 0 0.135514f
c54 4 0 0.00143442f
r55 70 74 0.660011
r56 47 56 1.16709
r57 47 74 11.3611
r58 42 70 2.37568
r59 39 42 1.16709
r60 32 56 0.0238214
r61 32 33 2.26917
r62 29 32 2.26917
r63 26 33 0.00605528
r64 24 29 0.00605528
r65 21 23 0.652036
r66 21 22 4.84305
r67 18 22 0.652036
r68 9 26 3.8511
r69 9 24 3.8511
r70 9 23 8.7525
r71 6 18 3.8511
r72 4 39 0.185659
r73 2 39 0.185659
.ends

.subckt PM_G4_XOR2_N2_B 2 4 7 10 19 20 28 31 35 45 52 55
c33 55 0 0.0280361f
c34 52 0 0.00155244f
c35 45 0 0.13326f
c36 35 0 0.154246f
c37 31 0 9.67975e-20
c38 28 0 0.117533f
c39 20 0 0.0348105f
c40 19 0 0.169544f
c41 10 0 0.209756f
c42 7 0 0.32787f
c43 4 0 0.134866f
c44 2 0 0.146861f
r45 49 55 1.16709
r46 49 52 0.0364688
r47 43 45 4.53833
r48 38 45 0.00605528
r49 35 47 1.87725
r50 33 47 0.527901
r51 32 43 0.00605528
r52 31 55 0.181909
r53 29 55 0.494161
r54 29 31 0.1167
r55 28 47 0.333556
r56 28 31 4.72635
r57 23 55 0.128424
r58 23 55 0.40845
r59 22 55 0.181909
r60 20 22 6.7686
r61 19 55 0.494161
r62 19 22 0.1167
r63 16 20 0.652036
r64 10 35 6.3018
r65 7 38 3.8511
r66 7 33 4.14285
r67 7 32 3.8511
r68 4 55 3.7344
r69 2 16 4.14285
.ends

.subckt PM_G4_XOR2_N2_Z 2 4 6 8 23 27 30 33
c29 30 0 0.00340522f
c30 27 0 0.00725263f
c31 23 0 0.0052085f
c32 8 0 0.00143442f
c33 6 0 0.00143442f
r34 33 35 3.83443
r35 30 33 6.00171
r36 27 35 1.16709
r37 23 30 1.16709
r38 8 27 0.185659
r39 6 23 0.185659
r40 4 27 0.185659
r41 2 23 0.185659
.ends

.subckt G4_XOR2_N2  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI14.X0 N_NET1_XI14.X0_D N_VDD_XI14.X0_PGD N_B_XI14.X0_CG N_VDD_XI14.X0_PGD
+ N_VSS_XI14.X0_S TIGFET_HPNW8
XI4.X0 N_NET2_XI4.X0_D N_VSS_XI4.X0_PGD N_A_XI4.X0_CG N_VSS_XI4.X0_PGD
+ N_VDD_XI4.X0_S TIGFET_HPNW8
XI12.X0 N_NET1_XI12.X0_D N_VSS_XI12.X0_PGD N_B_XI12.X0_CG N_VSS_XI12.X0_PGD
+ N_VDD_XI12.X0_S TIGFET_HPNW8
XI0.X0 N_NET2_XI0.X0_D N_VDD_XI0.X0_PGD N_A_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_B_XI15.X0_PGD N_NET2_XI15.X0_CG N_B_XI15.X0_PGD
+ N_VDD_XI15.X0_S TIGFET_HPNW8
XI6.X0 N_Z_XI6.X0_D N_A_XI6.X0_PGD N_B_XI6.X0_CG N_A_XI6.X0_PGD N_VSS_XI6.X0_S
+ TIGFET_HPNW8
XI13.X0 N_Z_XI13.X0_D N_NET1_XI13.X0_PGD N_A_XI13.X0_CG N_NET1_XI13.X0_PGD
+ N_VDD_XI13.X0_S TIGFET_HPNW8
XI2.X0 N_Z_XI2.X0_D N_NET2_XI2.X0_PGD N_NET1_XI2.X0_CG N_NET2_XI2.X0_PGD
+ N_VSS_XI2.X0_S TIGFET_HPNW8
*
x_PM_G4_XOR2_N2_VSS N_VSS_XI14.X0_S N_VSS_XI4.X0_PGD N_VSS_XI12.X0_PGD
+ N_VSS_XI0.X0_S N_VSS_XI6.X0_S N_VSS_XI2.X0_S N_VSS_c_5_p N_VSS_c_22_p
+ N_VSS_c_37_p N_VSS_c_4_p N_VSS_c_84_p N_VSS_c_7_p N_VSS_c_6_p N_VSS_c_91_p
+ N_VSS_c_8_p N_VSS_c_13_p N_VSS_c_29_p N_VSS_c_35_p N_VSS_c_39_p N_VSS_c_14_p
+ N_VSS_c_32_p N_VSS_c_9_p N_VSS_c_10_p N_VSS_c_18_p N_VSS_c_19_p N_VSS_c_25_p
+ N_VSS_c_28_p N_VSS_c_26_p N_VSS_c_55_p N_VSS_c_40_p N_VSS_c_77_p N_VSS_c_11_p
+ N_VSS_c_27_p VSS PM_G4_XOR2_N2_VSS
x_PM_G4_XOR2_N2_VDD N_VDD_XI14.X0_PGD N_VDD_XI4.X0_S N_VDD_XI12.X0_S
+ N_VDD_XI0.X0_PGD N_VDD_XI15.X0_S N_VDD_XI13.X0_S N_VDD_c_102_n N_VDD_c_149_p
+ N_VDD_c_103_n N_VDD_c_175_p N_VDD_c_104_n N_VDD_c_189_p N_VDD_c_105_n
+ N_VDD_c_110_n N_VDD_c_114_n N_VDD_c_117_n N_VDD_c_118_n N_VDD_c_119_n
+ N_VDD_c_126_n N_VDD_c_127_n N_VDD_c_128_n N_VDD_c_132_n N_VDD_c_135_n
+ N_VDD_c_154_p N_VDD_c_137_n N_VDD_c_162_p N_VDD_c_139_n N_VDD_c_140_n VDD
+ N_VDD_c_141_n N_VDD_c_143_n PM_G4_XOR2_N2_VDD
x_PM_G4_XOR2_N2_A N_A_XI4.X0_CG N_A_XI0.X0_CG N_A_XI6.X0_PGD N_A_XI13.X0_CG
+ N_A_c_198_n N_A_c_200_n N_A_c_201_n N_A_c_230_p N_A_c_216_n A N_A_c_202_n
+ N_A_c_204_n N_A_c_208_n N_A_c_209_n N_A_c_225_n N_A_c_229_p N_A_c_211_n
+ PM_G4_XOR2_N2_A
x_PM_G4_XOR2_N2_NET1 N_NET1_XI14.X0_D N_NET1_XI12.X0_D N_NET1_XI13.X0_PGD
+ N_NET1_XI2.X0_CG N_NET1_c_279_n N_NET1_c_263_n N_NET1_c_284_p N_NET1_c_256_n
+ N_NET1_c_257_n N_NET1_c_259_n N_NET1_c_273_n N_NET1_c_261_n PM_G4_XOR2_N2_NET1
x_PM_G4_XOR2_N2_NET2 N_NET2_XI4.X0_D N_NET2_XI0.X0_D N_NET2_XI15.X0_CG
+ N_NET2_XI2.X0_PGD N_NET2_c_315_n N_NET2_c_331_p N_NET2_c_316_n N_NET2_c_293_n
+ N_NET2_c_295_n N_NET2_c_299_n N_NET2_c_321_n N_NET2_c_303_n PM_G4_XOR2_N2_NET2
x_PM_G4_XOR2_N2_B N_B_XI14.X0_CG N_B_XI12.X0_CG N_B_XI15.X0_PGD N_B_XI6.X0_CG
+ N_B_c_338_n N_B_c_356_n N_B_c_340_n N_B_c_341_n N_B_c_358_n N_B_c_342_n B
+ N_B_c_345_n PM_G4_XOR2_N2_B
x_PM_G4_XOR2_N2_Z N_Z_XI15.X0_D N_Z_XI6.X0_D N_Z_XI13.X0_D N_Z_XI2.X0_D
+ N_Z_c_379_n N_Z_c_370_n N_Z_c_374_n Z PM_G4_XOR2_N2_Z
cc_1 N_VSS_XI4.X0_PGD N_VDD_XI14.X0_PGD 3.09777e-19
cc_2 N_VSS_XI12.X0_PGD N_VDD_XI14.X0_PGD 0.0019593f
cc_3 N_VSS_XI4.X0_PGD N_VDD_XI0.X0_PGD 0.0019696f
cc_4 N_VSS_c_4_p N_VDD_c_102_n 0.0019593f
cc_5 N_VSS_c_5_p N_VDD_c_103_n 0.0019696f
cc_6 N_VSS_c_6_p N_VDD_c_104_n 3.3848e-19
cc_7 N_VSS_c_7_p N_VDD_c_105_n 9.5668e-19
cc_8 N_VSS_c_8_p N_VDD_c_105_n 0.00165395f
cc_9 N_VSS_c_9_p N_VDD_c_105_n 0.00337557f
cc_10 N_VSS_c_10_p N_VDD_c_105_n 0.00738982f
cc_11 N_VSS_c_11_p N_VDD_c_105_n 9.16632e-19
cc_12 N_VSS_XI4.X0_PGD N_VDD_c_110_n 2.76462e-19
cc_13 N_VSS_c_13_p N_VDD_c_110_n 4.35319e-19
cc_14 N_VSS_c_14_p N_VDD_c_110_n 3.66936e-19
cc_15 N_VSS_c_10_p N_VDD_c_110_n 0.00312786f
cc_16 N_VSS_c_7_p N_VDD_c_114_n 3.4118e-19
cc_17 N_VSS_c_8_p N_VDD_c_114_n 4.19648e-19
cc_18 N_VSS_c_18_p N_VDD_c_114_n 0.0035394f
cc_19 N_VSS_c_19_p N_VDD_c_117_n 0.00106066f
cc_20 N_VSS_c_8_p N_VDD_c_118_n 5.20373e-19
cc_21 N_VSS_c_5_p N_VDD_c_119_n 3.9313e-19
cc_22 N_VSS_c_22_p N_VDD_c_119_n 3.9313e-19
cc_23 N_VSS_c_13_p N_VDD_c_119_n 0.00141228f
cc_24 N_VSS_c_14_p N_VDD_c_119_n 0.00114511f
cc_25 N_VSS_c_25_p N_VDD_c_119_n 0.00345257f
cc_26 N_VSS_c_26_p N_VDD_c_119_n 0.00601358f
cc_27 N_VSS_c_27_p N_VDD_c_119_n 7.74609e-19
cc_28 N_VSS_c_28_p N_VDD_c_126_n 0.00107662f
cc_29 N_VSS_c_29_p N_VDD_c_127_n 9.53862e-19
cc_30 N_VSS_c_4_p N_VDD_c_128_n 3.9313e-19
cc_31 N_VSS_c_29_p N_VDD_c_128_n 0.00161703f
cc_32 N_VSS_c_32_p N_VDD_c_128_n 2.26455e-19
cc_33 N_VSS_c_18_p N_VDD_c_128_n 0.0060445f
cc_34 N_VSS_c_13_p N_VDD_c_132_n 9.25722e-19
cc_35 N_VSS_c_35_p N_VDD_c_132_n 9.24903e-19
cc_36 N_VSS_c_14_p N_VDD_c_132_n 3.99794e-19
cc_37 N_VSS_c_37_p N_VDD_c_135_n 2.36788e-19
cc_38 N_VSS_c_29_p N_VDD_c_135_n 0.00251632f
cc_39 N_VSS_c_39_p N_VDD_c_137_n 2.22977e-19
cc_40 N_VSS_c_40_p N_VDD_c_137_n 0.00110879f
cc_41 N_VSS_c_10_p N_VDD_c_139_n 0.0010705f
cc_42 N_VSS_c_18_p N_VDD_c_140_n 0.00108916f
cc_43 N_VSS_c_29_p N_VDD_c_141_n 3.48267e-19
cc_44 N_VSS_c_32_p N_VDD_c_141_n 6.46219e-19
cc_45 N_VSS_c_13_p N_VDD_c_143_n 3.48267e-19
cc_46 N_VSS_c_14_p N_VDD_c_143_n 6.489e-19
cc_47 N_VSS_XI4.X0_PGD N_A_c_198_n 4.04227e-19
cc_48 N_VSS_XI12.X0_PGD N_A_c_198_n 2.49256e-19
cc_49 N_VSS_c_14_p N_A_c_200_n 9.46927e-19
cc_50 N_VSS_XI12.X0_PGD N_A_c_201_n 2.49256e-19
cc_51 N_VSS_c_13_p N_A_c_202_n 3.33636e-19
cc_52 N_VSS_c_14_p N_A_c_202_n 3.2351e-19
cc_53 N_VSS_c_35_p N_A_c_204_n 0.00580642f
cc_54 N_VSS_c_10_p N_A_c_204_n 7.28437e-19
cc_55 N_VSS_c_55_p N_A_c_204_n 0.00192457f
cc_56 N_VSS_c_40_p N_A_c_204_n 3.96468e-19
cc_57 N_VSS_c_55_p N_A_c_208_n 6.42713e-19
cc_58 N_VSS_c_13_p N_A_c_209_n 3.2351e-19
cc_59 N_VSS_c_14_p N_A_c_209_n 2.68747e-19
cc_60 N_VSS_c_55_p N_A_c_211_n 4.97622e-19
cc_61 N_VSS_c_7_p N_NET1_c_256_n 3.43419e-19
cc_62 N_VSS_c_8_p N_NET1_c_257_n 0.00115894f
cc_63 N_VSS_c_18_p N_NET1_c_257_n 2.79692e-19
cc_64 N_VSS_c_29_p N_NET1_c_259_n 0.00143375f
cc_65 N_VSS_c_35_p N_NET1_c_259_n 2.33463e-19
cc_66 N_VSS_c_9_p N_NET1_c_261_n 4.42442e-19
cc_67 N_VSS_c_18_p N_NET1_c_261_n 4.73555e-19
cc_68 N_VSS_c_6_p N_NET2_c_293_n 3.43419e-19
cc_69 N_VSS_c_35_p N_NET2_c_293_n 3.48267e-19
cc_70 N_VSS_c_6_p N_NET2_c_295_n 3.48267e-19
cc_71 N_VSS_c_35_p N_NET2_c_295_n 0.00163864f
cc_72 N_VSS_c_10_p N_NET2_c_295_n 6.00032e-19
cc_73 N_VSS_c_26_p N_NET2_c_295_n 2.79074e-19
cc_74 N_VSS_c_35_p N_NET2_c_299_n 0.00185959f
cc_75 N_VSS_c_26_p N_NET2_c_299_n 0.00111941f
cc_76 N_VSS_c_55_p N_NET2_c_299_n 0.0051115f
cc_77 N_VSS_c_77_p N_NET2_c_299_n 0.00115623f
cc_78 N_VSS_c_13_p N_NET2_c_303_n 5.67902e-19
cc_79 N_VSS_c_26_p N_NET2_c_303_n 4.76092e-19
cc_80 N_VSS_XI12.X0_PGD N_B_XI15.X0_PGD 0.00190378f
cc_81 N_VSS_XI4.X0_PGD N_B_c_338_n 2.59761e-19
cc_82 N_VSS_XI12.X0_PGD N_B_c_338_n 4.04459e-19
cc_83 N_VSS_XI12.X0_PGD N_B_c_340_n 4.08222e-19
cc_84 N_VSS_c_84_p N_B_c_341_n 8.74538e-19
cc_85 N_VSS_c_37_p N_B_c_342_n 0.00168656f
cc_86 N_VSS_c_29_p B 3.14335e-19
cc_87 N_VSS_c_32_p B 3.07907e-19
cc_88 N_VSS_c_29_p N_B_c_345_n 3.07907e-19
cc_89 N_VSS_c_32_p N_B_c_345_n 2.38856e-19
cc_90 N_VSS_c_6_p N_Z_c_370_n 3.43419e-19
cc_91 N_VSS_c_91_p N_Z_c_370_n 3.43419e-19
cc_92 N_VSS_c_35_p N_Z_c_370_n 3.48267e-19
cc_93 N_VSS_c_39_p N_Z_c_370_n 3.48267e-19
cc_94 N_VSS_c_6_p N_Z_c_374_n 3.48267e-19
cc_95 N_VSS_c_91_p N_Z_c_374_n 3.48267e-19
cc_96 N_VSS_c_35_p N_Z_c_374_n 4.84964e-19
cc_97 N_VSS_c_39_p N_Z_c_374_n 5.71987e-19
cc_98 N_VSS_c_55_p N_Z_c_374_n 3.24575e-19
cc_99 N_VDD_XI0.X0_PGD N_A_XI6.X0_PGD 0.00170367f
cc_100 N_VDD_XI14.X0_PGD N_A_c_198_n 2.49256e-19
cc_101 N_VDD_XI0.X0_PGD N_A_c_198_n 4.07423e-19
cc_102 N_VDD_XI0.X0_PGD N_A_c_201_n 4.08222e-19
cc_103 N_VDD_c_149_p N_A_c_216_n 0.00170367f
cc_104 N_VDD_c_105_n N_A_c_202_n 5.04211e-19
cc_105 N_VDD_c_127_n N_A_c_202_n 2.0061e-19
cc_106 N_VDD_c_132_n N_A_c_204_n 4.55539e-19
cc_107 N_VDD_c_143_n N_A_c_204_n 3.5189e-19
cc_108 N_VDD_c_154_p N_A_c_208_n 6.92642e-19
cc_109 N_VDD_c_105_n N_A_c_209_n 5.74039e-19
cc_110 N_VDD_c_127_n N_A_c_209_n 2.00694e-19
cc_111 N_VDD_c_141_n N_A_c_209_n 2.58157e-19
cc_112 N_VDD_c_132_n N_A_c_225_n 4.08069e-19
cc_113 N_VDD_c_143_n N_A_c_225_n 6.61916e-19
cc_114 N_VDD_c_154_p N_A_c_211_n 8.87092e-19
cc_115 N_VDD_c_154_p N_NET1_c_263_n 8.59992e-19
cc_116 N_VDD_c_162_p N_NET1_c_263_n 2.76493e-19
cc_117 N_VDD_c_104_n N_NET1_c_256_n 3.43419e-19
cc_118 N_VDD_c_135_n N_NET1_c_256_n 3.48267e-19
cc_119 N_VDD_c_104_n N_NET1_c_257_n 3.48267e-19
cc_120 N_VDD_c_128_n N_NET1_c_257_n 4.34701e-19
cc_121 N_VDD_c_135_n N_NET1_c_257_n 0.00119216f
cc_122 N_VDD_c_135_n N_NET1_c_259_n 0.00121188f
cc_123 N_VDD_c_154_p N_NET1_c_259_n 0.00357992f
cc_124 N_VDD_c_162_p N_NET1_c_259_n 8.17443e-19
cc_125 N_VDD_c_135_n N_NET1_c_273_n 2.78343e-19
cc_126 N_VDD_c_154_p N_NET1_c_273_n 2.67643e-19
cc_127 N_VDD_c_162_p N_NET1_c_273_n 3.70842e-19
cc_128 N_VDD_c_127_n N_NET1_c_261_n 2.94681e-19
cc_129 N_VDD_c_175_p N_NET2_c_293_n 3.67949e-19
cc_130 N_VDD_c_118_n N_NET2_c_293_n 3.72199e-19
cc_131 N_VDD_c_175_p N_NET2_c_295_n 3.9802e-19
cc_132 N_VDD_c_118_n N_NET2_c_295_n 5.226e-19
cc_133 N_VDD_c_119_n N_NET2_c_295_n 4.34701e-19
cc_134 N_VDD_c_132_n N_NET2_c_299_n 2.89449e-19
cc_135 N_VDD_c_105_n N_B_XI14.X0_CG 3.86879e-19
cc_136 N_VDD_XI14.X0_PGD N_B_c_338_n 4.0747e-19
cc_137 N_VDD_XI0.X0_PGD N_B_c_338_n 2.59761e-19
cc_138 N_VDD_XI0.X0_PGD N_B_c_340_n 2.59761e-19
cc_139 N_VDD_c_135_n N_B_c_342_n 2.45557e-19
cc_140 N_VDD_c_154_p N_B_c_342_n 0.00104936f
cc_141 N_VDD_c_143_n N_B_c_345_n 3.88194e-19
cc_142 N_VDD_c_104_n N_Z_c_379_n 3.43419e-19
cc_143 N_VDD_c_189_p N_Z_c_379_n 3.43419e-19
cc_144 N_VDD_c_135_n N_Z_c_379_n 3.48267e-19
cc_145 N_VDD_c_154_p N_Z_c_379_n 3.4118e-19
cc_146 N_VDD_c_137_n N_Z_c_379_n 3.72199e-19
cc_147 N_VDD_c_104_n N_Z_c_374_n 3.48267e-19
cc_148 N_VDD_c_189_p N_Z_c_374_n 3.48267e-19
cc_149 N_VDD_c_135_n N_Z_c_374_n 7.9714e-19
cc_150 N_VDD_c_154_p N_Z_c_374_n 6.28755e-19
cc_151 N_VDD_c_137_n N_Z_c_374_n 8.5731e-19
cc_152 N_A_XI13.X0_CG N_NET1_XI13.X0_PGD 9.16948e-19
cc_153 N_A_c_229_p N_NET1_XI13.X0_PGD 5.82245e-19
cc_154 N_A_c_230_p N_NET1_c_279_n 8.72031e-19
cc_155 N_A_c_208_n N_NET1_c_259_n 0.00253116f
cc_156 N_A_c_211_n N_NET1_c_259_n 6.96104e-19
cc_157 N_A_c_229_p N_NET1_c_273_n 2.38856e-19
cc_158 N_A_XI13.X0_CG N_NET2_XI15.X0_CG 2.29068e-19
cc_159 N_A_XI6.X0_PGD N_NET2_XI2.X0_PGD 0.00174971f
cc_160 N_A_c_201_n N_NET2_XI2.X0_PGD 3.14428e-19
cc_161 N_A_c_229_p N_NET2_XI2.X0_PGD 3.71891e-19
cc_162 N_A_XI6.X0_PGD N_NET2_c_315_n 4.63684e-19
cc_163 N_A_c_216_n N_NET2_c_316_n 0.00174971f
cc_164 N_A_c_198_n N_NET2_c_293_n 5.99889e-19
cc_165 N_A_c_204_n N_NET2_c_299_n 0.0021219f
cc_166 N_A_c_208_n N_NET2_c_299_n 0.00109012f
cc_167 N_A_c_225_n N_NET2_c_299_n 3.44698e-19
cc_168 N_A_c_230_p N_NET2_c_321_n 4.27572e-19
cc_169 N_A_c_204_n N_NET2_c_321_n 3.44698e-19
cc_170 N_A_c_225_n N_NET2_c_321_n 6.78604e-19
cc_171 N_A_c_201_n N_B_XI6.X0_CG 0.003858f
cc_172 N_A_c_198_n N_B_c_338_n 0.00631299f
cc_173 N_A_c_209_n N_B_c_356_n 8.20069e-19
cc_174 N_A_c_201_n N_B_c_340_n 0.00464284f
cc_175 N_A_c_201_n N_B_c_358_n 0.00220484f
cc_176 N_A_c_198_n N_B_c_345_n 8.92181e-19
cc_177 N_A_c_204_n N_Z_c_374_n 0.00336431f
cc_178 N_A_c_208_n N_Z_c_374_n 0.00291096f
cc_179 N_A_c_229_p N_Z_c_374_n 9.75659e-19
cc_180 N_NET1_XI13.X0_PGD N_NET2_XI15.X0_CG 2.3921e-19
cc_181 N_NET1_c_284_p N_NET2_XI2.X0_PGD 0.00790765f
cc_182 N_NET1_XI13.X0_PGD N_NET2_c_315_n 0.00383f
cc_183 N_NET1_c_256_n N_NET2_c_293_n 2.51993e-19
cc_184 N_NET1_XI13.X0_PGD N_B_XI15.X0_PGD 0.00215865f
cc_185 N_NET1_XI2.X0_CG N_B_XI6.X0_CG 2.58346e-19
cc_186 N_NET1_c_256_n N_B_c_338_n 5.53604e-19
cc_187 N_NET1_c_284_p N_B_c_358_n 2.58346e-19
cc_188 N_NET1_c_263_n N_B_c_342_n 0.00193302f
cc_189 N_NET1_c_259_n N_Z_c_374_n 2.36895e-19
cc_190 N_NET2_XI15.X0_CG N_B_XI15.X0_PGD 0.00204226f
cc_191 N_NET2_c_315_n N_B_XI15.X0_PGD 0.00161654f
cc_192 N_NET2_XI2.X0_PGD N_B_c_358_n 0.00351134f
cc_193 N_NET2_c_331_p N_B_c_358_n 0.00396313f
cc_194 N_NET2_c_315_n N_Z_c_379_n 7.46018e-19
cc_195 N_NET2_c_315_n N_Z_c_370_n 2.51166e-19
cc_196 N_NET2_XI2.X0_PGD N_Z_c_374_n 0.0012102f
cc_197 N_NET2_c_315_n N_Z_c_374_n 2.5304e-19
cc_198 N_NET2_c_299_n N_Z_c_374_n 3.59687e-19
cc_199 N_B_c_358_n N_Z_c_374_n 0.00106974f
*
.ends
*
*
.subckt XOR2_HPNW8 A B Y VDD VSS
xgate (VSS VDD A B Y) G4_XOR2_N2
.ends
*
* File: G5_XOR3_N2.pex.netlist
* Created: Thu Mar 31 11:38:36 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XOR3_N2_VDD 2 5 9 12 14 17 34 35 44 45 47 54 55 65 69 74 77 79 80
+ 81 84 86 90 93 96 98 102 104 108 112 114 116 118 119 125 134 139 Vss
c115 139 Vss 0.00504502f
c116 134 Vss 0.00507145f
c117 125 Vss 0.00564924f
c118 119 Vss 2.39889e-19
c119 118 Vss 4.91626e-19
c120 117 Vss 5.50975e-19
c121 114 Vss 4.52364e-19
c122 112 Vss 0.00169191f
c123 108 Vss 0.00106552f
c124 104 Vss 0.00630988f
c125 102 Vss 0.00113412f
c126 98 Vss 0.00579331f
c127 96 Vss 0.00150773f
c128 93 Vss 0.00256047f
c129 90 Vss 0.00487749f
c130 86 Vss 0.00657827f
c131 84 Vss 0.00152345f
c132 81 Vss 8.67722e-19
c133 80 Vss 0.00905163f
c134 79 Vss 0.0103203f
c135 77 Vss 0.00223293f
c136 74 Vss 0.00377995f
c137 69 Vss 0.00394389f
c138 65 Vss 0.00382792f
c139 55 Vss 0.035607f
c140 54 Vss 0.100823f
c141 47 Vss 8.75732e-20
c142 45 Vss 0.0356105f
c143 44 Vss 0.101295f
c144 35 Vss 0.0346386f
c145 34 Vss 0.0990802f
c146 17 Vss 0.269219f
c147 9 Vss 0.270254f
c148 5 Vss 0.27424f
r149 110 112 5.2515
r150 108 139 1.16709
r151 106 108 2.16729
r152 105 119 0.494161
r153 104 110 0.652036
r154 104 105 7.46046
r155 102 134 1.16709
r156 100 119 0.128424
r157 100 102 2.16729
r158 99 118 0.494161
r159 98 106 0.652036
r160 98 99 10.3363
r161 94 117 0.0828784
r162 94 96 2.00578
r163 93 118 0.128424
r164 92 117 0.551426
r165 92 93 4.58464
r166 90 125 1.16709
r167 88 117 0.551426
r168 88 90 6.79361
r169 87 116 0.326018
r170 86 118 0.494161
r171 86 87 10.1279
r172 82 114 0.0828784
r173 82 84 1.82344
r174 80 119 0.494161
r175 80 81 15.8795
r176 79 116 0.326018
r177 78 114 0.551426
r178 78 79 15.6295
r179 77 114 0.551426
r180 76 81 0.652036
r181 76 77 4.58464
r182 74 112 1.16709
r183 69 96 1.16709
r184 65 84 1.16709
r185 57 139 0.0476429
r186 55 57 1.45875
r187 54 58 0.652036
r188 54 57 1.45875
r189 51 55 0.652036
r190 47 134 0.0476429
r191 45 47 1.45875
r192 44 48 0.652036
r193 44 47 1.45875
r194 41 45 0.652036
r195 37 125 0.238214
r196 35 37 1.45875
r197 34 38 0.652036
r198 34 37 1.45875
r199 31 35 0.652036
r200 17 58 3.8511
r201 17 51 3.8511
r202 14 74 0.185659
r203 12 69 0.185659
r204 9 48 3.8511
r205 9 41 3.8511
r206 5 38 3.8511
r207 5 31 3.8511
r208 2 65 0.185659
.ends

.subckt PM_G5_XOR3_N2_C 2 4 6 8 17 20 23 32 37 40 43 47 52 57 84 92 98 Vss
c55 98 Vss 3.07681e-19
c56 92 Vss 0.00543335f
c57 84 Vss 0.00807877f
c58 57 Vss 0.00478462f
c59 52 Vss 0.00202371f
c60 47 Vss 0.00149319f
c61 43 Vss 5.64514e-19
c62 40 Vss 6.40888e-19
c63 37 Vss 0.00399277f
c64 32 Vss 0.00492048f
c65 23 Vss 2.41681e-19
c66 20 Vss 0.221837f
c67 17 Vss 0.126125f
c68 15 Vss 0.0247918f
c69 4 Vss 0.133869f
r70 93 98 0.441572
r71 92 94 0.655813
r72 92 93 9.04425
r73 88 98 0.174814
r74 84 98 0.441572
r75 52 94 2.45904
r76 47 88 2.45904
r77 43 57 1.16709
r78 43 84 22.1365
r79 40 43 0.0416786
r80 37 52 1.16709
r81 32 47 1.16709
r82 23 57 0.0476429
r83 21 23 0.326018
r84 21 23 0.1167
r85 20 24 0.652036
r86 20 23 6.7686
r87 17 57 0.357321
r88 15 23 0.326018
r89 15 17 0.40845
r90 8 37 0.185659
r91 6 32 0.185659
r92 4 24 3.8511
r93 2 17 3.44265
.ends

.subckt PM_G5_XOR3_N2_VSS 3 6 8 11 15 18 34 37 44 45 54 55 57 66 70 73 78 83 88
+ 93 98 107 112 121 123 124 125 130 131 136 142 148 152 153 154 156 Vss
c125 154 Vss 3.75522e-19
c126 153 Vss 3.88979e-19
c127 152 Vss 4.4306e-19
c128 148 Vss 4.18562e-19
c129 142 Vss 0.00192878f
c130 136 Vss 0.00349848f
c131 131 Vss 8.4146e-19
c132 130 Vss 0.00631713f
c133 125 Vss 8.38522e-19
c134 124 Vss 0.00567123f
c135 123 Vss 0.00379369f
c136 121 Vss 0.00292495f
c137 112 Vss 0.00392167f
c138 107 Vss 0.00408825f
c139 98 Vss 0.00496033f
c140 93 Vss 0.00183916f
c141 88 Vss 6.78589e-19
c142 83 Vss 8.07476e-19
c143 78 Vss 0.00294517f
c144 73 Vss 0.00293431f
c145 70 Vss 0.00527641f
c146 66 Vss 0.00738472f
c147 57 Vss 1.05421e-19
c148 55 Vss 0.0347733f
c149 54 Vss 0.0996929f
c150 45 Vss 0.035088f
c151 44 Vss 0.0994129f
c152 37 Vss 6.29003e-20
c153 35 Vss 0.0348882f
c154 34 Vss 0.100326f
c155 15 Vss 0.270318f
c156 11 Vss 0.269056f
c157 8 Vss 0.00143442f
c158 3 Vss 0.275257f
r159 148 156 0.326018
r160 143 154 0.494161
r161 142 156 0.326018
r162 142 143 7.46046
r163 138 154 0.128424
r164 137 153 0.494161
r165 136 144 0.652036
r166 136 137 7.46046
r167 132 153 0.128424
r168 130 154 0.494161
r169 130 131 15.8795
r170 126 152 0.0828784
r171 124 153 0.494161
r172 124 125 13.0037
r173 123 131 0.652036
r174 122 152 0.551426
r175 122 123 12.0451
r176 121 152 0.551426
r177 120 125 0.652036
r178 120 121 8.169
r179 93 148 5.2515
r180 88 112 1.16709
r181 88 144 2.16729
r182 83 107 1.16709
r183 83 138 2.16729
r184 78 132 5.2515
r185 73 98 1.16709
r186 73 126 4.33978
r187 70 93 1.16709
r188 66 78 1.16709
r189 57 112 0.0476429
r190 55 57 1.45875
r191 54 58 0.652036
r192 54 57 1.45875
r193 51 55 0.652036
r194 47 107 0.0476429
r195 45 47 1.45875
r196 44 48 0.652036
r197 44 47 1.45875
r198 41 45 0.652036
r199 37 98 0.238214
r200 35 37 1.45875
r201 34 38 0.652036
r202 34 37 1.45875
r203 31 35 0.652036
r204 18 70 0.185659
r205 15 58 3.8511
r206 15 51 3.8511
r207 11 48 3.8511
r208 11 41 3.8511
r209 8 66 0.185659
r210 6 66 0.185659
r211 3 38 3.8511
r212 3 31 3.8511
.ends

.subckt PM_G5_XOR3_N2_CI 2 4 6 8 23 26 31 34 39 44 79 80 82 84 89 Vss
c55 95 Vss 8.69704e-20
c56 89 Vss 0.00497463f
c57 84 Vss 1.28221e-19
c58 83 Vss 1.74838e-19
c59 82 Vss 0.0011265f
c60 80 Vss 4.20409e-19
c61 79 Vss 0.00494114f
c62 44 Vss 0.00209131f
c63 39 Vss 0.00145787f
c64 34 Vss 0.00360912f
c65 31 Vss 0.00501643f
c66 26 Vss 0.00386883f
c67 23 Vss 0.00546777f
c68 4 Vss 0.00143442f
r69 90 95 0.494161
r70 89 91 0.652036
r71 89 90 10.3363
r72 85 95 0.128424
r73 83 95 0.494161
r74 83 84 1.70882
r75 82 84 0.652036
r76 81 82 4.75136
r77 79 81 0.652036
r78 79 80 18.9638
r79 75 80 0.652036
r80 44 91 2.58407
r81 39 85 2.58407
r82 34 75 7.71054
r83 31 44 1.16709
r84 26 39 1.16709
r85 23 34 1.16709
r86 8 31 0.185659
r87 6 26 0.185659
r88 4 23 0.185659
r89 2 23 0.185659
.ends

.subckt PM_G5_XOR3_N2_A 2 4 7 11 24 44 45 49 51 54 56 57 60 65 66 69 74 Vss
c72 74 Vss 0.00550397f
c73 69 Vss 0.00508271f
c74 66 Vss 0.00601821f
c75 65 Vss 3.90863e-19
c76 57 Vss 9.08254e-19
c77 56 Vss 6.01198e-19
c78 54 Vss 0.00400006f
c79 51 Vss 0.00786937f
c80 49 Vss 0.135055f
c81 45 Vss 0.127825f
c82 44 Vss 9.84889e-20
c83 24 Vss 0.21954f
c84 21 Vss 0.129208f
c85 19 Vss 0.0247918f
c86 7 Vss 1.22248f
c87 4 Vss 0.139574f
r88 65 74 1.16709
r89 65 66 0.531835
r90 62 69 1.16709
r91 60 62 0.0416786
r92 57 60 0.833571
r93 56 66 10.4613
r94 53 56 0.652036
r95 53 54 8.66914
r96 52 57 0.0685365
r97 51 54 0.652036
r98 51 52 10.2113
r99 47 49 4.53833
r100 44 74 0.0238214
r101 44 45 2.26917
r102 41 44 2.26917
r103 36 49 0.00605528
r104 35 45 0.00605528
r105 32 47 0.00605528
r106 31 41 0.00605528
r107 27 69 0.0952857
r108 25 27 0.326018
r109 25 27 0.1167
r110 24 28 0.652036
r111 24 27 6.7686
r112 21 27 0.3335
r113 19 27 0.326018
r114 19 21 0.2334
r115 11 36 3.8511
r116 11 32 3.8511
r117 7 11 15.4044
r118 7 35 3.8511
r119 7 11 15.4044
r120 7 31 3.8511
r121 4 28 3.8511
r122 2 21 3.6177
.ends

.subckt PM_G5_XOR3_N2_BI 2 4 6 8 18 21 29 32 37 42 51 56 65 71 72 80 Vss
c67 80 Vss 3.59704e-19
c68 72 Vss 1.29652e-19
c69 71 Vss 7.91966e-19
c70 65 Vss 0.00113976f
c71 56 Vss 0.00255458f
c72 51 Vss 0.00236417f
c73 42 Vss 0.00116078f
c74 37 Vss 0.00223673f
c75 32 Vss 0.00202587f
c76 29 Vss 0.00450527f
c77 21 Vss 0.111942f
c78 6 Vss 0.112114f
c79 4 Vss 0.00143442f
r80 76 80 0.655813
r81 71 72 0.655813
r82 70 71 3.501
r83 65 70 0.655813
r84 42 56 1.16709
r85 42 72 2.00578
r86 37 51 1.16709
r87 37 80 12.0712
r88 37 65 2.00578
r89 32 76 2.45904
r90 29 32 1.16709
r91 21 56 0.50025
r92 18 51 0.50025
r93 8 21 3.09255
r94 6 18 3.09255
r95 4 29 0.185659
r96 2 29 0.185659
.ends

.subckt PM_G5_XOR3_N2_AI 2 4 7 11 31 37 43 46 51 60 73 79 Vss
c46 79 Vss 2.59226e-19
c47 73 Vss 0.00489127f
c48 60 Vss 0.00532163f
c49 51 Vss 0.00226804f
c50 46 Vss 0.00262268f
c51 43 Vss 0.00448639f
c52 37 Vss 0.127877f
c53 31 Vss 0.131547f
c54 7 Vss 1.20882f
c55 4 Vss 0.00143442f
r56 75 79 0.652036
r57 73 79 13.7539
r58 51 60 1.16709
r59 51 73 2.75079
r60 46 75 5.2515
r61 43 46 1.16709
r62 36 60 0.0238214
r63 36 37 2.334
r64 33 36 2.20433
r65 29 31 4.53833
r66 26 37 0.00605528
r67 25 31 0.00605528
r68 22 33 0.00605528
r69 21 29 0.00605528
r70 11 26 3.8511
r71 11 22 3.8511
r72 7 11 15.4044
r73 7 25 3.8511
r74 7 11 15.4044
r75 7 21 3.8511
r76 4 43 0.185659
r77 2 43 0.185659
.ends

.subckt PM_G5_XOR3_N2_B 2 4 6 8 16 17 24 26 33 38 42 45 50 55 60 65 73 74 80 86
+ 91 92 Vss
c75 92 Vss 1.50842e-19
c76 91 Vss 6.9543e-19
c77 86 Vss 8.71217e-19
c78 80 Vss 6.55917e-19
c79 74 Vss 5.2356e-19
c80 73 Vss 0.00528129f
c81 65 Vss 0.00250661f
c82 60 Vss 0.00217314f
c83 55 Vss 0.00427742f
c84 50 Vss 0.00149379f
c85 45 Vss 3.19996e-19
c86 42 Vss 4.98048e-19
c87 38 Vss 6.6601e-19
c88 33 Vss 1.05421e-19
c89 26 Vss 0.111942f
c90 24 Vss 9.84889e-20
c91 20 Vss 0.0247918f
c92 17 Vss 0.0339811f
c93 16 Vss 0.183683f
c94 8 Vss 0.111942f
c95 4 Vss 0.12597f
c96 2 Vss 0.136912f
r97 90 92 0.655813
r98 90 91 3.501
r99 86 91 0.655813
r100 73 80 0.0685365
r101 73 74 10.3363
r102 69 74 0.652036
r103 50 65 1.16709
r104 50 92 2.00578
r105 45 60 1.16709
r106 45 86 2.00578
r107 45 80 2.04225
r108 38 55 1.16709
r109 38 69 2.25064
r110 38 42 0.0364688
r111 36 55 0.0476429
r112 33 65 0.50025
r113 26 60 0.50025
r114 24 55 0.357321
r115 20 36 0.326018
r116 20 24 0.40845
r117 17 36 6.7686
r118 16 36 0.326018
r119 16 36 0.1167
r120 13 17 0.652036
r121 8 33 3.09255
r122 6 26 3.09255
r123 4 24 3.44265
r124 2 13 3.8511
.ends

.subckt PM_G5_XOR3_N2_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00368262f
c33 27 Vss 0.00842339f
c34 23 Vss 0.00745376f
c35 8 Vss 0.00143442f
c36 6 Vss 0.00334862f
r37 33 35 5.20982
r38 30 40 1.16709
r39 30 33 5.79332
r40 27 35 1.16709
r41 23 40 0.05
r42 8 27 0.185659
r43 6 23 0.185659
r44 4 27 0.185659
r45 2 23 0.185659
.ends

.subckt G5_XOR3_N2  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI15.X0 N_CI_XI15.X0_D N_VSS_XI15.X0_PGD N_C_XI15.X0_CG N_VSS_XI15.X0_PGD
+ N_VDD_XI15.X0_S TIGFET_HPNW8
XI12.X0 N_CI_XI12.X0_D N_VDD_XI12.X0_PGD N_C_XI12.X0_CG N_VDD_XI12.X0_PGD
+ N_VSS_XI12.X0_S TIGFET_HPNW8
XI11.X0 N_BI_XI11.X0_D N_VDD_XI11.X0_PGD N_B_XI11.X0_CG N_VDD_XI11.X0_PGD
+ N_VSS_XI11.X0_S TIGFET_HPNW8
XI13.X0 N_AI_XI13.X0_D N_VSS_XI13.X0_PGD N_A_XI13.X0_CG N_VSS_XI13.X0_PGD
+ N_VDD_XI13.X0_S TIGFET_HPNW8
XI14.X0 N_BI_XI14.X0_D N_VSS_XI14.X0_PGD N_B_XI14.X0_CG N_VSS_XI14.X0_PGD
+ N_VDD_XI14.X0_S TIGFET_HPNW8
XI0.X0 N_AI_XI0.X0_D N_VDD_XI0.X0_PGD N_A_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW8
XI18.X0 N_Z_XI18.X0_D N_AI_XI18.X0_PGD N_BI_XI18.X0_CG N_AI_XI18.X0_PGD
+ N_C_XI18.X0_S TIGFET_HPNW8
XI16.X0 N_Z_XI16.X0_D N_AI_XI16.X0_PGD N_B_XI16.X0_CG N_AI_XI16.X0_PGD
+ N_CI_XI16.X0_S TIGFET_HPNW8
XI19.X0 N_Z_XI19.X0_D N_A_XI19.X0_PGD N_B_XI19.X0_CG N_A_XI19.X0_PGD
+ N_C_XI19.X0_S TIGFET_HPNW8
XI17.X0 N_Z_XI17.X0_D N_A_XI17.X0_PGD N_BI_XI17.X0_CG N_A_XI17.X0_PGD
+ N_CI_XI17.X0_S TIGFET_HPNW8
*
x_PM_G5_XOR3_N2_VDD N_VDD_XI15.X0_S N_VDD_XI12.X0_PGD N_VDD_XI11.X0_PGD
+ N_VDD_XI13.X0_S N_VDD_XI14.X0_S N_VDD_XI0.X0_PGD N_VDD_c_112_p N_VDD_c_20_p
+ N_VDD_c_25_p N_VDD_c_4_p N_VDD_c_93_p N_VDD_c_102_p N_VDD_c_21_p N_VDD_c_75_p
+ N_VDD_c_103_p N_VDD_c_6_p N_VDD_c_7_p N_VDD_c_13_p N_VDD_c_5_p N_VDD_c_62_p
+ N_VDD_c_30_p N_VDD_c_63_p N_VDD_c_31_p N_VDD_c_17_p N_VDD_c_64_p N_VDD_c_22_p
+ N_VDD_c_10_p N_VDD_c_26_p N_VDD_c_38_p N_VDD_c_11_p N_VDD_c_58_p VDD
+ N_VDD_c_66_p N_VDD_c_70_p N_VDD_c_2_p N_VDD_c_43_p N_VDD_c_39_p Vss
+ PM_G5_XOR3_N2_VDD
x_PM_G5_XOR3_N2_C N_C_XI15.X0_CG N_C_XI12.X0_CG N_C_XI18.X0_S N_C_XI19.X0_S
+ N_C_c_134_p N_C_c_118_n N_C_c_128_p N_C_c_121_n N_C_c_165_p C N_C_c_130_p
+ N_C_c_148_p N_C_c_167_p N_C_c_124_n N_C_c_125_n N_C_c_150_p N_C_c_154_p Vss
+ PM_G5_XOR3_N2_C
x_PM_G5_XOR3_N2_VSS N_VSS_XI15.X0_PGD N_VSS_XI12.X0_S N_VSS_XI11.X0_S
+ N_VSS_XI13.X0_PGD N_VSS_XI14.X0_PGD N_VSS_XI0.X0_S N_VSS_c_179_n N_VSS_c_235_n
+ N_VSS_c_180_n N_VSS_c_182_n N_VSS_c_183_n N_VSS_c_184_n N_VSS_c_289_p
+ N_VSS_c_186_n N_VSS_c_252_p N_VSS_c_187_n N_VSS_c_192_n N_VSS_c_195_n
+ N_VSS_c_199_n N_VSS_c_203_n N_VSS_c_204_n N_VSS_c_207_n N_VSS_c_211_n
+ N_VSS_c_215_n N_VSS_c_218_n N_VSS_c_220_n N_VSS_c_221_n N_VSS_c_222_n
+ N_VSS_c_226_n N_VSS_c_227_n N_VSS_c_230_n N_VSS_c_286_p N_VSS_c_231_n
+ N_VSS_c_232_n N_VSS_c_233_n VSS Vss PM_G5_XOR3_N2_VSS
x_PM_G5_XOR3_N2_CI N_CI_XI15.X0_D N_CI_XI12.X0_D N_CI_XI16.X0_S N_CI_XI17.X0_S
+ N_CI_c_296_n N_CI_c_309_n N_CI_c_343_p N_CI_c_298_n N_CI_c_316_n N_CI_c_345_p
+ N_CI_c_302_n N_CI_c_319_n N_CI_c_320_n N_CI_c_333_p N_CI_c_326_p Vss
+ PM_G5_XOR3_N2_CI
x_PM_G5_XOR3_N2_A N_A_XI13.X0_CG N_A_XI0.X0_CG N_A_XI19.X0_PGD N_A_XI17.X0_PGD
+ N_A_c_351_n N_A_c_405_p N_A_c_396_p N_A_c_398_p N_A_c_352_n N_A_c_358_n
+ N_A_c_359_n N_A_c_360_n A N_A_c_367_n N_A_c_368_n N_A_c_361_n N_A_c_410_p Vss
+ PM_G5_XOR3_N2_A
x_PM_G5_XOR3_N2_BI N_BI_XI11.X0_D N_BI_XI14.X0_D N_BI_XI18.X0_CG N_BI_XI17.X0_CG
+ N_BI_c_446_n N_BI_c_447_n N_BI_c_423_n N_BI_c_426_n N_BI_c_430_n N_BI_c_443_n
+ N_BI_c_453_n N_BI_c_455_n N_BI_c_433_n N_BI_c_476_p N_BI_c_444_n N_BI_c_434_n
+ Vss PM_G5_XOR3_N2_BI
x_PM_G5_XOR3_N2_AI N_AI_XI13.X0_D N_AI_XI0.X0_D N_AI_XI18.X0_PGD
+ N_AI_XI16.X0_PGD N_AI_c_500_n N_AI_c_491_n N_AI_c_492_n N_AI_c_494_n
+ N_AI_c_507_n N_AI_c_530_p N_AI_c_498_n N_AI_c_510_n Vss PM_G5_XOR3_N2_AI
x_PM_G5_XOR3_N2_B N_B_XI11.X0_CG N_B_XI14.X0_CG N_B_XI16.X0_CG N_B_XI19.X0_CG
+ N_B_c_537_n N_B_c_538_n N_B_c_546_n N_B_c_600_n N_B_c_564_n N_B_c_539_n B
+ N_B_c_580_n N_B_c_554_n N_B_c_540_n N_B_c_585_n N_B_c_572_n N_B_c_541_n
+ N_B_c_556_n N_B_c_557_n N_B_c_543_n N_B_c_597_n N_B_c_544_n Vss
+ PM_G5_XOR3_N2_B
x_PM_G5_XOR3_N2_Z N_Z_XI18.X0_D N_Z_XI16.X0_D N_Z_XI19.X0_D N_Z_XI17.X0_D
+ N_Z_c_611_n N_Z_c_618_n N_Z_c_615_n Z Vss PM_G5_XOR3_N2_Z
cc_1 N_VDD_XI11.X0_PGD N_C_XI12.X0_CG 0.00111653f
cc_2 N_VDD_c_2_p N_C_XI12.X0_CG 9.52277e-19
cc_3 N_VDD_XI12.X0_PGD N_C_c_118_n 4.18724e-19
cc_4 N_VDD_c_4_p N_C_c_118_n 0.00111653f
cc_5 N_VDD_c_5_p N_C_c_118_n 0.00134893f
cc_6 N_VDD_c_6_p N_C_c_121_n 3.43419e-19
cc_7 N_VDD_c_7_p C 4.76491e-19
cc_8 N_VDD_c_5_p C 0.00161703f
cc_9 N_VDD_c_5_p N_C_c_124_n 2.84956e-19
cc_10 N_VDD_c_10_p N_C_c_125_n 4.83409e-19
cc_11 N_VDD_c_11_p N_C_c_125_n 7.93016e-19
cc_12 N_VDD_XI12.X0_PGD N_VSS_XI15.X0_PGD 0.00201307f
cc_13 N_VDD_c_13_p N_VSS_XI15.X0_PGD 3.1461e-19
cc_14 N_VDD_c_5_p N_VSS_XI15.X0_PGD 2.01827e-19
cc_15 N_VDD_XI11.X0_PGD N_VSS_XI13.X0_PGD 2.35243e-19
cc_16 N_VDD_XI0.X0_PGD N_VSS_XI13.X0_PGD 0.00201252f
cc_17 N_VDD_c_17_p N_VSS_XI13.X0_PGD 3.00522e-19
cc_18 N_VDD_XI11.X0_PGD N_VSS_XI14.X0_PGD 0.00200584f
cc_19 N_VDD_XI0.X0_PGD N_VSS_XI14.X0_PGD 2.22638e-19
cc_20 N_VDD_c_20_p N_VSS_c_179_n 0.00201307f
cc_21 N_VDD_c_21_p N_VSS_c_180_n 0.00201252f
cc_22 N_VDD_c_22_p N_VSS_c_180_n 2.84671e-19
cc_23 N_VDD_c_22_p N_VSS_c_182_n 3.9313e-19
cc_24 N_VDD_c_11_p N_VSS_c_183_n 2.41035e-19
cc_25 N_VDD_c_25_p N_VSS_c_184_n 0.00200584f
cc_26 N_VDD_c_26_p N_VSS_c_184_n 3.9313e-19
cc_27 N_VDD_c_5_p N_VSS_c_186_n 3.4118e-19
cc_28 N_VDD_c_13_p N_VSS_c_187_n 4.32468e-19
cc_29 N_VDD_c_5_p N_VSS_c_187_n 3.85027e-19
cc_30 N_VDD_c_30_p N_VSS_c_187_n 0.00120518f
cc_31 N_VDD_c_31_p N_VSS_c_187_n 3.98949e-19
cc_32 N_VDD_c_2_p N_VSS_c_187_n 3.48267e-19
cc_33 N_VDD_c_5_p N_VSS_c_192_n 3.98099e-19
cc_34 N_VDD_c_10_p N_VSS_c_192_n 7.43603e-19
cc_35 N_VDD_c_11_p N_VSS_c_192_n 5.11768e-19
cc_36 N_VDD_c_17_p N_VSS_c_195_n 6.74818e-19
cc_37 N_VDD_c_22_p N_VSS_c_195_n 0.00161703f
cc_38 N_VDD_c_38_p N_VSS_c_195_n 8.6926e-19
cc_39 N_VDD_c_39_p N_VSS_c_195_n 3.48267e-19
cc_40 N_VDD_c_10_p N_VSS_c_199_n 6.78479e-19
cc_41 N_VDD_c_26_p N_VSS_c_199_n 0.00161703f
cc_42 N_VDD_c_11_p N_VSS_c_199_n 0.00242479f
cc_43 N_VDD_c_43_p N_VSS_c_199_n 3.48267e-19
cc_44 N_VDD_c_38_p N_VSS_c_203_n 7.32365e-19
cc_45 N_VDD_c_13_p N_VSS_c_204_n 4.41003e-19
cc_46 N_VDD_c_31_p N_VSS_c_204_n 3.89161e-19
cc_47 N_VDD_c_2_p N_VSS_c_204_n 7.99831e-19
cc_48 N_VDD_c_17_p N_VSS_c_207_n 3.48267e-19
cc_49 N_VDD_c_22_p N_VSS_c_207_n 2.26455e-19
cc_50 N_VDD_c_38_p N_VSS_c_207_n 3.99794e-19
cc_51 N_VDD_c_39_p N_VSS_c_207_n 6.489e-19
cc_52 N_VDD_c_10_p N_VSS_c_211_n 3.82294e-19
cc_53 N_VDD_c_26_p N_VSS_c_211_n 2.26455e-19
cc_54 N_VDD_c_11_p N_VSS_c_211_n 9.55109e-19
cc_55 N_VDD_c_43_p N_VSS_c_211_n 6.46219e-19
cc_56 N_VDD_c_7_p N_VSS_c_215_n 0.00347459f
cc_57 N_VDD_c_13_p N_VSS_c_215_n 0.00229697f
cc_58 N_VDD_c_58_p N_VSS_c_215_n 0.0010705f
cc_59 N_VDD_c_13_p N_VSS_c_218_n 0.0086177f
cc_60 N_VDD_c_31_p N_VSS_c_218_n 0.00116809f
cc_61 N_VDD_c_5_p N_VSS_c_220_n 0.00954271f
cc_62 N_VDD_c_62_p N_VSS_c_221_n 0.00107367f
cc_63 N_VDD_c_63_p N_VSS_c_222_n 0.00827847f
cc_64 N_VDD_c_64_p N_VSS_c_222_n 7.30484e-19
cc_65 N_VDD_c_22_p N_VSS_c_222_n 0.00369102f
cc_66 N_VDD_c_66_p N_VSS_c_222_n 0.00149929f
cc_67 N_VDD_c_13_p N_VSS_c_226_n 0.0010758f
cc_68 N_VDD_c_5_p N_VSS_c_227_n 0.00143208f
cc_69 N_VDD_c_26_p N_VSS_c_227_n 0.00601868f
cc_70 N_VDD_c_70_p N_VSS_c_227_n 0.00107091f
cc_71 N_VDD_c_22_p N_VSS_c_230_n 0.00534674f
cc_72 N_VDD_c_13_p N_VSS_c_231_n 0.00112682f
cc_73 N_VDD_c_5_p N_VSS_c_232_n 0.00107375f
cc_74 N_VDD_c_22_p N_VSS_c_233_n 7.74609e-19
cc_75 N_VDD_c_75_p N_CI_c_296_n 3.43419e-19
cc_76 N_VDD_c_30_p N_CI_c_296_n 3.72199e-19
cc_77 N_VDD_c_75_p N_CI_c_298_n 3.48267e-19
cc_78 N_VDD_c_5_p N_CI_c_298_n 4.34701e-19
cc_79 N_VDD_c_30_p N_CI_c_298_n 5.226e-19
cc_80 N_VDD_c_31_p N_CI_c_298_n 0.00101464f
cc_81 N_VDD_c_31_p N_CI_c_302_n 6.82638e-19
cc_82 N_VDD_c_64_p N_CI_c_302_n 7.0762e-19
cc_83 N_VDD_XI0.X0_PGD N_A_c_351_n 3.94784e-19
cc_84 N_VDD_XI0.X0_PGD N_A_c_352_n 2.73656e-19
cc_85 N_VDD_c_6_p N_A_c_352_n 2.69869e-19
cc_86 N_VDD_c_22_p N_A_c_352_n 4.57714e-19
cc_87 N_VDD_c_38_p N_A_c_352_n 3.99109e-19
cc_88 N_VDD_c_11_p N_A_c_352_n 3.90005e-19
cc_89 N_VDD_c_39_p N_A_c_352_n 2.43883e-19
cc_90 N_VDD_c_6_p N_A_c_358_n 9.18655e-19
cc_91 N_VDD_c_11_p N_A_c_359_n 0.00564482f
cc_92 N_VDD_c_31_p N_A_c_360_n 0.00104501f
cc_93 N_VDD_c_93_p N_A_c_361_n 3.61944e-19
cc_94 N_VDD_c_31_p N_A_c_361_n 5.71421e-19
cc_95 N_VDD_c_6_p N_BI_c_423_n 3.43419e-19
cc_96 N_VDD_c_26_p N_BI_c_423_n 3.4118e-19
cc_97 N_VDD_c_11_p N_BI_c_423_n 3.48267e-19
cc_98 N_VDD_c_6_p N_BI_c_426_n 3.48267e-19
cc_99 N_VDD_c_26_p N_BI_c_426_n 3.98099e-19
cc_100 N_VDD_c_11_p N_BI_c_426_n 4.99861e-19
cc_101 N_VDD_XI0.X0_PGD N_AI_XI18.X0_PGD 3.2392e-19
cc_102 N_VDD_c_102_p N_AI_c_491_n 3.2392e-19
cc_103 N_VDD_c_103_p N_AI_c_492_n 3.43419e-19
cc_104 N_VDD_c_64_p N_AI_c_492_n 3.73302e-19
cc_105 N_VDD_c_103_p N_AI_c_494_n 3.48267e-19
cc_106 N_VDD_c_64_p N_AI_c_494_n 5.23123e-19
cc_107 N_VDD_c_22_p N_AI_c_494_n 4.34701e-19
cc_108 N_VDD_c_38_p N_AI_c_494_n 5.44192e-19
cc_109 N_VDD_c_22_p N_AI_c_498_n 4.11874e-19
cc_110 N_VDD_XI12.X0_PGD N_B_XI11.X0_CG 0.00111821f
cc_111 N_VDD_XI11.X0_PGD N_B_c_537_n 3.99339e-19
cc_112 N_VDD_c_112_p N_B_c_538_n 0.00111821f
cc_113 N_VDD_c_31_p N_B_c_539_n 7.52847e-19
cc_114 N_VDD_c_39_p N_B_c_540_n 4.92948e-19
cc_115 N_VDD_c_11_p N_B_c_541_n 3.15013e-19
cc_116 N_C_c_118_n N_VSS_XI15.X0_PGD 4.18724e-19
cc_117 N_C_c_128_p N_VSS_c_235_n 4.96533e-19
cc_118 C N_VSS_c_187_n 2.70019e-19
cc_119 N_C_c_130_p N_VSS_c_187_n 2.56587e-19
cc_120 N_C_c_125_n N_VSS_c_187_n 2.07529e-19
cc_121 N_C_c_125_n N_VSS_c_192_n 0.00194391f
cc_122 N_C_c_125_n N_VSS_c_199_n 0.00158941f
cc_123 N_C_c_134_p N_VSS_c_204_n 0.00249737f
cc_124 C N_VSS_c_204_n 2.87758e-19
cc_125 N_C_c_124_n N_VSS_c_204_n 2.0363e-19
cc_126 N_C_c_130_p N_VSS_c_215_n 4.01014e-19
cc_127 N_C_c_125_n N_VSS_c_215_n 2.67374e-19
cc_128 C N_VSS_c_220_n 3.52403e-19
cc_129 N_C_c_130_p N_VSS_c_220_n 0.00136475f
cc_130 N_C_c_125_n N_VSS_c_220_n 0.00317947f
cc_131 N_C_c_125_n N_VSS_c_227_n 0.00191592f
cc_132 N_C_c_118_n N_CI_c_296_n 6.55689e-19
cc_133 N_C_c_125_n N_CI_c_298_n 0.00101026f
cc_134 N_C_c_125_n N_CI_c_302_n 0.00289054f
cc_135 N_C_c_125_n N_A_c_352_n 2.24413e-19
cc_136 N_C_c_121_n N_A_c_358_n 8.20481e-19
cc_137 N_C_c_148_p N_A_c_358_n 0.00195474f
cc_138 N_C_c_125_n N_A_c_359_n 4.776e-19
cc_139 N_C_c_150_p N_A_c_367_n 2.7748e-19
cc_140 N_C_c_148_p N_A_c_368_n 0.0018313f
cc_141 N_C_c_125_n N_A_c_368_n 3.28319e-19
cc_142 N_C_c_150_p N_A_c_368_n 0.00220096f
cc_143 N_C_c_154_p N_A_c_368_n 2.81326e-19
cc_144 N_C_c_125_n N_BI_c_426_n 0.00113193f
cc_145 N_C_c_148_p N_BI_c_430_n 0.00119554f
cc_146 N_C_c_125_n N_BI_c_430_n 0.00400118f
cc_147 N_C_c_150_p N_BI_c_430_n 6.70289e-19
cc_148 N_C_c_150_p N_BI_c_433_n 8.45766e-19
cc_149 N_C_c_125_n N_BI_c_434_n 6.63379e-19
cc_150 N_C_c_148_p N_B_c_541_n 4.44753e-19
cc_151 N_C_c_150_p N_B_c_543_n 3.99616e-19
cc_152 N_C_c_150_p N_B_c_544_n 0.00180761f
cc_153 N_C_c_121_n N_Z_c_611_n 3.43419e-19
cc_154 N_C_c_165_p N_Z_c_611_n 3.43419e-19
cc_155 N_C_c_148_p N_Z_c_611_n 3.48267e-19
cc_156 N_C_c_167_p N_Z_c_611_n 3.48267e-19
cc_157 N_C_c_165_p N_Z_c_615_n 3.48267e-19
cc_158 N_C_c_148_p N_Z_c_615_n 6.09821e-19
cc_159 N_C_c_167_p N_Z_c_615_n 5.71987e-19
cc_160 N_VSS_c_186_n N_CI_c_296_n 3.43419e-19
cc_161 N_VSS_c_192_n N_CI_c_296_n 3.48267e-19
cc_162 N_VSS_c_252_p N_CI_c_309_n 3.43419e-19
cc_163 N_VSS_c_186_n N_CI_c_298_n 3.48267e-19
cc_164 N_VSS_c_187_n N_CI_c_298_n 5.88914e-19
cc_165 N_VSS_c_192_n N_CI_c_298_n 8.10527e-19
cc_166 N_VSS_c_215_n N_CI_c_298_n 4.71364e-19
cc_167 N_VSS_c_218_n N_CI_c_298_n 9.66309e-19
cc_168 N_VSS_c_220_n N_CI_c_298_n 2.82247e-19
cc_169 N_VSS_c_203_n N_CI_c_316_n 8.74405e-19
cc_170 N_VSS_c_195_n N_CI_c_302_n 3.79792e-19
cc_171 N_VSS_c_230_n N_CI_c_302_n 5.41979e-19
cc_172 N_VSS_c_222_n N_CI_c_319_n 0.00182487f
cc_173 N_VSS_c_203_n N_CI_c_320_n 0.00142004f
cc_174 N_VSS_XI13.X0_PGD N_A_c_351_n 3.91587e-19
cc_175 N_VSS_c_203_n N_A_c_352_n 8.4508e-19
cc_176 N_VSS_c_230_n N_A_c_352_n 4.69076e-19
cc_177 N_VSS_c_195_n N_A_c_360_n 3.32273e-19
cc_178 N_VSS_c_207_n N_A_c_360_n 3.1261e-19
cc_179 N_VSS_c_195_n N_A_c_361_n 3.04912e-19
cc_180 N_VSS_c_207_n N_A_c_361_n 0.00110478f
cc_181 N_VSS_c_186_n N_BI_c_423_n 3.43419e-19
cc_182 N_VSS_c_192_n N_BI_c_423_n 3.48267e-19
cc_183 N_VSS_c_186_n N_BI_c_426_n 3.48267e-19
cc_184 N_VSS_c_192_n N_BI_c_426_n 8.10527e-19
cc_185 N_VSS_c_227_n N_BI_c_426_n 2.79692e-19
cc_186 N_VSS_XI14.X0_PGD N_AI_XI18.X0_PGD 2.74627e-19
cc_187 N_VSS_c_183_n N_AI_c_500_n 2.74627e-19
cc_188 N_VSS_c_252_p N_AI_c_492_n 3.43419e-19
cc_189 N_VSS_c_203_n N_AI_c_492_n 3.48267e-19
cc_190 N_VSS_c_252_p N_AI_c_494_n 3.48267e-19
cc_191 N_VSS_c_195_n N_AI_c_494_n 0.00108072f
cc_192 N_VSS_c_203_n N_AI_c_494_n 0.00213737f
cc_193 N_VSS_c_230_n N_AI_c_494_n 2.86662e-19
cc_194 N_VSS_c_203_n N_AI_c_507_n 0.00122373f
cc_195 N_VSS_c_230_n N_AI_c_498_n 0.00370204f
cc_196 N_VSS_c_286_p N_AI_c_498_n 0.0017148f
cc_197 N_VSS_c_230_n N_AI_c_510_n 0.0018958f
cc_198 N_VSS_XI14.X0_PGD N_B_c_537_n 3.96142e-19
cc_199 N_VSS_c_289_p N_B_c_546_n 9.56171e-19
cc_200 N_VSS_c_199_n N_B_c_539_n 2.57202e-19
cc_201 N_VSS_c_199_n B 3.42746e-19
cc_202 N_VSS_c_211_n B 3.2351e-19
cc_203 N_VSS_c_199_n N_B_c_540_n 3.2351e-19
cc_204 N_VSS_c_211_n N_B_c_540_n 2.68747e-19
cc_205 N_VSS_c_203_n N_B_c_541_n 3.58501e-19
cc_206 N_CI_c_302_n N_A_c_352_n 0.00183351f
cc_207 N_CI_c_302_n N_A_c_360_n 3.36095e-19
cc_208 N_CI_c_298_n N_BI_c_426_n 9.23808e-19
cc_209 N_CI_c_316_n N_BI_c_430_n 2.81279e-19
cc_210 N_CI_c_302_n N_BI_c_430_n 0.0032559f
cc_211 N_CI_c_326_p N_BI_c_443_n 8.83269e-19
cc_212 N_CI_c_326_p N_BI_c_444_n 2.18743e-19
cc_213 N_CI_c_302_n N_BI_c_434_n 0.00153557f
cc_214 N_CI_c_302_n N_AI_c_494_n 0.00135858f
cc_215 N_CI_c_320_n N_AI_c_494_n 0.00128778f
cc_216 N_CI_c_326_p N_AI_c_507_n 0.00144463f
cc_217 N_CI_c_302_n N_AI_c_498_n 0.00198979f
cc_218 N_CI_c_333_p N_AI_c_498_n 0.00533258f
cc_219 N_CI_c_326_p N_AI_c_498_n 0.00290048f
cc_220 N_CI_c_298_n N_B_c_539_n 5.51453e-19
cc_221 N_CI_c_326_p N_B_c_554_n 6.37546e-19
cc_222 N_CI_c_316_n N_B_c_541_n 5.58533e-19
cc_223 N_CI_c_302_n N_B_c_556_n 0.00108926f
cc_224 N_CI_c_326_p N_B_c_557_n 2.05643e-19
cc_225 N_CI_c_302_n N_B_c_543_n 4.54861e-19
cc_226 N_CI_c_326_p N_B_c_543_n 0.00179506f
cc_227 N_CI_c_309_n N_Z_c_618_n 3.43419e-19
cc_228 N_CI_c_343_p N_Z_c_618_n 3.43419e-19
cc_229 N_CI_c_316_n N_Z_c_618_n 3.48267e-19
cc_230 N_CI_c_345_p N_Z_c_618_n 3.48267e-19
cc_231 N_CI_c_309_n N_Z_c_615_n 3.48267e-19
cc_232 N_CI_c_343_p N_Z_c_615_n 3.48267e-19
cc_233 N_CI_c_316_n N_Z_c_615_n 5.71987e-19
cc_234 N_CI_c_345_p N_Z_c_615_n 5.71987e-19
cc_235 N_CI_c_302_n N_Z_c_615_n 4.15391e-19
cc_236 N_A_c_368_n N_BI_c_446_n 2.74063e-19
cc_237 N_A_XI19.X0_PGD N_BI_c_447_n 9.65637e-19
cc_238 N_A_c_352_n N_BI_c_426_n 3.85685e-19
cc_239 N_A_c_358_n N_BI_c_426_n 4.22951e-19
cc_240 N_A_c_358_n N_BI_c_430_n 0.00110458f
cc_241 N_A_c_368_n N_BI_c_430_n 8.05288e-19
cc_242 N_A_c_368_n N_BI_c_443_n 2.98812e-19
cc_243 N_A_c_358_n N_BI_c_453_n 3.37713e-19
cc_244 N_A_c_368_n N_BI_c_453_n 2.96819e-19
cc_245 N_A_XI19.X0_PGD N_BI_c_455_n 0.00133285f
cc_246 N_A_c_368_n N_BI_c_433_n 0.00102169f
cc_247 N_A_c_352_n N_BI_c_434_n 4.10091e-19
cc_248 N_A_XI19.X0_PGD N_AI_XI18.X0_PGD 0.0174244f
cc_249 N_A_c_358_n N_AI_XI18.X0_PGD 9.55469e-19
cc_250 N_A_c_368_n N_AI_XI18.X0_PGD 7.53964e-19
cc_251 N_A_c_396_p N_AI_c_500_n 0.00199315f
cc_252 N_A_c_368_n N_AI_c_500_n 0.00125772f
cc_253 N_A_c_398_p N_AI_c_491_n 0.00201004f
cc_254 N_A_c_351_n N_AI_c_492_n 6.89066e-19
cc_255 N_A_c_352_n N_AI_c_494_n 7.80381e-19
cc_256 N_A_XI19.X0_PGD N_B_XI19.X0_CG 9.65637e-19
cc_257 N_A_c_351_n N_B_c_537_n 0.0035308f
cc_258 N_A_c_352_n N_B_c_537_n 6.06747e-19
cc_259 N_A_c_361_n N_B_c_538_n 5.83549e-19
cc_260 N_A_c_405_p N_B_c_564_n 9.37683e-19
cc_261 N_A_c_358_n N_B_c_539_n 6.35249e-19
cc_262 N_A_c_352_n B 9.05205e-19
cc_263 N_A_c_358_n B 5.05926e-19
cc_264 N_A_c_367_n N_B_c_554_n 5.53953e-19
cc_265 N_A_c_410_p N_B_c_554_n 3.2351e-19
cc_266 N_A_c_351_n N_B_c_540_n 9.10729e-19
cc_267 N_A_c_358_n N_B_c_540_n 6.84646e-19
cc_268 N_A_XI19.X0_PGD N_B_c_572_n 0.00133285f
cc_269 N_A_c_410_p N_B_c_572_n 2.68747e-19
cc_270 N_A_c_352_n N_B_c_541_n 0.00336092f
cc_271 N_A_c_358_n N_B_c_541_n 0.00192865f
cc_272 N_A_c_368_n N_B_c_541_n 8.22275e-19
cc_273 N_A_c_352_n N_B_c_556_n 5.17628e-19
cc_274 N_A_c_368_n N_Z_c_611_n 0.00107687f
cc_275 N_A_XI19.X0_PGD N_Z_c_615_n 7.94638e-19
cc_276 N_A_c_358_n N_Z_c_615_n 0.00143807f
cc_277 N_A_c_368_n N_Z_c_615_n 0.0014359f
cc_278 N_BI_XI18.X0_CG N_AI_XI18.X0_PGD 9.47088e-19
cc_279 N_BI_c_453_n N_AI_XI18.X0_PGD 0.00133285f
cc_280 N_BI_c_430_n N_AI_c_498_n 9.24953e-19
cc_281 N_BI_c_423_n N_B_c_537_n 6.89066e-19
cc_282 N_BI_c_430_n N_B_c_539_n 0.00155724f
cc_283 N_BI_c_430_n N_B_c_580_n 6.02887e-19
cc_284 N_BI_c_444_n N_B_c_580_n 3.08318e-19
cc_285 N_BI_c_443_n N_B_c_554_n 0.0017864f
cc_286 N_BI_c_455_n N_B_c_554_n 4.56568e-19
cc_287 N_BI_c_433_n N_B_c_554_n 0.00165721f
cc_288 N_BI_c_430_n N_B_c_585_n 4.56568e-19
cc_289 N_BI_c_453_n N_B_c_585_n 0.00266356f
cc_290 N_BI_c_455_n N_B_c_585_n 7.16621e-19
cc_291 N_BI_c_453_n N_B_c_572_n 6.17967e-19
cc_292 N_BI_c_455_n N_B_c_572_n 0.00243716f
cc_293 N_BI_c_430_n N_B_c_541_n 0.00391901f
cc_294 N_BI_c_430_n N_B_c_557_n 3.07174e-19
cc_295 N_BI_c_433_n N_B_c_557_n 0.00126004f
cc_296 N_BI_c_476_p N_B_c_557_n 0.00342237f
cc_297 N_BI_c_430_n N_B_c_543_n 5.09978e-19
cc_298 N_BI_c_433_n N_B_c_543_n 7.34826e-19
cc_299 N_BI_c_444_n N_B_c_543_n 8.56575e-19
cc_300 N_BI_c_476_p N_B_c_597_n 0.00210118f
cc_301 N_BI_c_430_n N_B_c_544_n 0.00142766f
cc_302 N_BI_c_433_n N_B_c_544_n 9.32988e-19
cc_303 N_BI_c_430_n N_Z_c_615_n 0.00138952f
cc_304 N_BI_c_443_n N_Z_c_615_n 0.00138952f
cc_305 N_BI_c_453_n N_Z_c_615_n 8.66889e-19
cc_306 N_BI_c_455_n N_Z_c_615_n 8.66889e-19
cc_307 N_BI_c_433_n N_Z_c_615_n 0.00103509f
cc_308 N_BI_c_476_p N_Z_c_615_n 0.00212989f
cc_309 N_BI_c_444_n N_Z_c_615_n 0.00103331f
cc_310 N_AI_XI18.X0_PGD N_B_c_600_n 9.65637e-19
cc_311 N_AI_c_507_n N_B_c_580_n 3.6769e-19
cc_312 N_AI_c_530_p N_B_c_580_n 3.2351e-19
cc_313 N_AI_XI18.X0_PGD N_B_c_585_n 0.00133285f
cc_314 N_AI_c_507_n N_B_c_585_n 3.2351e-19
cc_315 N_AI_c_530_p N_B_c_585_n 0.00117301f
cc_316 N_AI_c_507_n N_B_c_557_n 4.82497e-19
cc_317 N_AI_XI18.X0_PGD N_Z_c_615_n 4.32017e-19
cc_318 N_B_c_580_n N_Z_c_615_n 0.00157325f
cc_319 N_B_c_554_n N_Z_c_615_n 0.00138952f
cc_320 N_B_c_572_n N_Z_c_615_n 8.66889e-19
cc_321 N_B_c_557_n N_Z_c_615_n 4.69528e-19
*
.ends
*
*
.subckt XOR3_HPNW8 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XOR3_N2
.ends
