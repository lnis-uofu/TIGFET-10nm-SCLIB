* sclib_tigfet10_hpall_tt_0p70v_25c.sp
.subckt TIGFET_HPNW1 D PGD CG PGS S
xgate (D PGD CG PGS S) TIGFET nw=1
.ends
.subckt TIGFET_HPNW4 D PGD CG PGS S
xgate (D PGD CG PGS S) TIGFET nw=4
.ends
.subckt TIGFET_HPNW8 D PGD CG PGS S
xgate (D PGD CG PGS S) TIGFET nw=8
.ends
.subckt TIGFET_HPNW12 D PGD CG PGS S
xgate (D PGD CG PGS S) TIGFET nw=12
.ends
*
* File: G3_AND2_N1.pex.netlist
* Created: Wed Feb 23 10:37:48 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_AND2_N1_VSS 2 4 6 8 10 12 14 16 30 31 33 50 53 70 75 80 85 94 99
+ 108 109 113 114 119 125 127 132 133 134 136 Vss
c68 134 Vss 3.75522e-19
c69 133 Vss 3.62111e-19
c70 132 Vss 0.00361417f
c71 127 Vss 0.00255728f
c72 125 Vss 0.00548072f
c73 119 Vss 0.00398592f
c74 114 Vss 9.65205e-19
c75 113 Vss 0.00179171f
c76 109 Vss 8.2274e-19
c77 108 Vss 0.00426189f
c78 99 Vss 0.00393602f
c79 94 Vss 0.004332f
c80 85 Vss 7.10513e-22
c81 80 Vss 6.65776e-19
c82 75 Vss 3.89225e-19
c83 70 Vss 0.00133027f
c84 58 Vss 0.0299355f
c85 57 Vss 0.0299355f
c86 53 Vss 7.50699e-20
c87 51 Vss 0.0346861f
c88 50 Vss 0.0984533f
c89 42 Vss 0.105926f
c90 37 Vss 0.0688517f
c91 33 Vss 6.52493e-20
c92 31 Vss 0.0342473f
c93 30 Vss 0.064644f
c94 16 Vss 0.00266844f
c95 14 Vss 0.0828881f
c96 12 Vss 0.0825199f
c97 10 Vss 0.0830027f
c98 8 Vss 0.0831275f
c99 6 Vss 0.0832632f
c100 4 Vss 0.0828837f
c101 2 Vss 0.00266829f
r102 132 136 0.326018
r103 131 132 4.16786
r104 127 131 0.655813
r105 126 134 0.494161
r106 125 136 0.326018
r107 125 126 10.1279
r108 121 134 0.128424
r109 120 133 0.494161
r110 119 134 0.494161
r111 119 120 10.378
r112 115 133 0.128424
r113 113 133 0.494161
r114 113 114 4.37625
r115 108 114 0.668428
r116 107 109 0.6565
r117 107 108 10.093
r118 85 127 1.82344
r119 80 99 1.16709
r120 80 121 2.16729
r121 75 94 1.16709
r122 75 115 2.16729
r123 70 109 1.85991
r124 53 99 0.238214
r125 51 53 1.45875
r126 50 54 0.652036
r127 50 53 1.45875
r128 47 51 0.652036
r129 43 58 0.494161
r130 42 44 0.652036
r131 42 43 2.9175
r132 39 58 0.128424
r133 38 57 0.494161
r134 37 58 0.494161
r135 37 38 2.8008
r136 34 57 0.128424
r137 33 94 0.238214
r138 31 33 1.4004
r139 30 57 0.494161
r140 30 33 1.5171
r141 27 31 0.652036
r142 16 85 1.16709
r143 14 47 2.5674
r144 12 54 2.5674
r145 10 44 2.5674
r146 8 39 2.5674
r147 6 27 2.5674
r148 4 34 2.5674
r149 2 70 1.16709
.ends

.subckt PM_G3_AND2_N1_VDD 2 4 6 10 12 25 27 33 51 53 54 58 60 64 68 70 74 76 78
+ 79 85 94 Vss
c87 94 Vss 0.00555165f
c88 85 Vss 0.00507125f
c89 79 Vss 4.42156e-19
c90 76 Vss 5.947e-19
c91 74 Vss 0.00125165f
c92 70 Vss 0.00410186f
c93 68 Vss 0.0014864f
c94 64 Vss 0.0023623f
c95 60 Vss 0.00679469f
c96 58 Vss 0.0016182f
c97 55 Vss 0.00207011f
c98 54 Vss 0.0101277f
c99 53 Vss 0.0036687f
c100 51 Vss 0.00587536f
c101 33 Vss 0.0347789f
c102 32 Vss 0.101192f
c103 27 Vss 0.183894f
c104 25 Vss 0.0364084f
c105 12 Vss 0.0842982f
c106 10 Vss 0.0825186f
c107 6 Vss 0.00153036f
c108 4 Vss 0.00221866f
c109 2 Vss 0.0976708f
r110 74 94 1.16709
r111 72 74 2.16729
r112 71 79 0.494161
r113 70 72 0.652036
r114 70 71 7.46046
r115 66 79 0.128424
r116 66 68 4.83471
r117 64 85 1.16709
r118 62 64 3.66771
r119 61 78 0.386734
r120 60 79 0.494161
r121 60 61 13.0037
r122 56 76 0.18826
r123 56 58 1.82344
r124 54 62 0.652036
r125 54 55 10.0862
r126 53 78 0.284962
r127 52 76 0.427332
r128 52 53 3.07105
r129 51 76 0.427332
r130 50 55 0.671696
r131 50 51 7.86189
r132 35 94 0.238214
r133 33 35 1.45875
r134 32 36 0.652036
r135 32 35 1.45875
r136 29 33 0.652036
r137 27 85 0.50025
r138 25 27 5.11257
r139 22 25 0.652541
r140 12 36 2.5674
r141 10 29 2.5674
r142 6 68 1.16709
r143 4 58 1.16709
r144 2 22 3.2676
.ends

.subckt PM_G3_AND2_N1_A 2 4 10 13 18 21 26 31 Vss
c25 31 Vss 0.00351715f
c26 26 Vss 0.00299969f
c27 18 Vss 8.55683e-19
c28 13 Vss 0.0576606f
c29 2 Vss 0.0575116f
r30 23 31 1.16709
r31 21 23 2.12561
r32 18 26 1.16709
r33 18 21 2.70911
r34 13 31 0.50025
r35 10 26 0.50025
r36 4 13 1.80885
r37 2 10 1.80885
.ends

.subckt PM_G3_AND2_N1_NET1 2 4 8 10 21 24 27 45 53 66 70 Vss
c51 70 Vss 0.00676771f
c52 66 Vss 0.00607266f
c53 53 Vss 0.00254578f
c54 45 Vss 0.00159242f
c55 27 Vss 1.04894e-19
c56 24 Vss 0.225594f
c57 21 Vss 0.0713786f
c58 19 Vss 0.0247918f
c59 10 Vss 0.0847975f
c60 4 Vss 0.00148239f
c61 2 Vss 0.00144265f
r62 70 74 0.652036
r63 53 66 1.16709
r64 53 74 3.66771
r65 48 70 8.04396
r66 48 50 6.4185
r67 45 48 2.75079
r68 27 66 0.0476429
r69 25 27 0.326018
r70 25 27 0.1167
r71 24 28 0.652036
r72 24 27 6.7686
r73 21 66 0.357321
r74 19 27 0.326018
r75 19 21 0.40845
r76 10 28 2.5674
r77 8 21 2.15895
r78 4 50 1.16709
r79 2 45 1.16709
.ends

.subckt PM_G3_AND2_N1_B 2 4 10 11 14 18 21 Vss
c26 21 Vss 5.0923e-19
c27 14 Vss 0.148163f
c28 11 Vss 0.0348321f
c29 10 Vss 0.287297f
c30 2 Vss 0.172263f
r31 18 21 0.0364688
r32 14 21 1.16709
r33 12 14 2.8008
r34 10 12 0.652036
r35 10 11 8.92755
r36 7 11 0.652036
r37 4 14 3.0342
r38 2 7 5.835
.ends

.subckt PM_G3_AND2_N1_Z 2 16 19 Vss
c11 2 Vss 0.00148239f
r12 16 19 0.0364688
r13 2 19 1.16709
.ends

.subckt G3_AND2_N1  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI7.X0 N_NET1_XI7.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_B_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW1
XI8.X0 N_NET1_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW1
XI9.X0 N_NET1_XI8.X0_D N_VSS_XI9.X0_PGD N_B_XI9.X0_CG N_VSS_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW1
XI2.X0 N_Z_XI2.X0_D N_VSS_XI2.X0_PGD N_NET1_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW1
XI1.X0 N_Z_XI2.X0_D N_VDD_XI1.X0_PGD N_NET1_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
*
x_PM_G3_AND2_N1_VSS N_VSS_XI7.X0_S N_VSS_XI8.X0_PGD N_VSS_XI8.X0_PGS
+ N_VSS_XI9.X0_PGD N_VSS_XI9.X0_PGS N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI1.X0_S N_VSS_c_13_p N_VSS_c_14_p N_VSS_c_42_p N_VSS_c_2_p N_VSS_c_49_p
+ N_VSS_c_4_p N_VSS_c_7_p N_VSS_c_23_p N_VSS_c_65_p N_VSS_c_8_p N_VSS_c_25_p
+ N_VSS_c_5_p N_VSS_c_6_p N_VSS_c_17_p N_VSS_c_10_p N_VSS_c_18_p N_VSS_c_30_p
+ N_VSS_c_68_p N_VSS_c_33_p N_VSS_c_19_p N_VSS_c_31_p VSS Vss PM_G3_AND2_N1_VSS
x_PM_G3_AND2_N1_VDD N_VDD_XI7.X0_PGD N_VDD_XI8.X0_S N_VDD_XI9.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_c_143_p N_VDD_c_128_p N_VDD_c_70_n
+ N_VDD_c_71_n N_VDD_c_75_n N_VDD_c_79_n N_VDD_c_80_n N_VDD_c_81_n N_VDD_c_116_p
+ N_VDD_c_88_n N_VDD_c_94_n N_VDD_c_100_n N_VDD_c_102_n VDD N_VDD_c_103_n
+ N_VDD_c_113_p N_VDD_c_104_n Vss PM_G3_AND2_N1_VDD
x_PM_G3_AND2_N1_A N_A_XI7.X0_CG N_A_XI8.X0_CG N_A_c_164_n N_A_c_156_n
+ N_A_c_157_n A N_A_c_167_n N_A_c_160_n Vss PM_G3_AND2_N1_A
x_PM_G3_AND2_N1_NET1 N_NET1_XI7.X0_D N_NET1_XI8.X0_D N_NET1_XI2.X0_CG
+ N_NET1_XI1.X0_CG N_NET1_c_183_n N_NET1_c_184_n N_NET1_c_185_n N_NET1_c_187_n
+ N_NET1_c_190_n N_NET1_c_193_n N_NET1_c_195_n Vss PM_G3_AND2_N1_NET1
x_PM_G3_AND2_N1_B N_B_XI7.X0_PGS N_B_XI9.X0_CG N_B_c_232_n N_B_c_234_n
+ N_B_c_239_n B N_B_c_242_n Vss PM_G3_AND2_N1_B
x_PM_G3_AND2_N1_Z N_Z_XI2.X0_D Z N_Z_c_260_n Vss PM_G3_AND2_N1_Z
cc_1 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.0016786f
cc_2 N_VSS_c_2_p N_VDD_c_70_n 0.0016786f
cc_3 N_VSS_XI7.X0_S N_VDD_c_71_n 9.73142e-19
cc_4 N_VSS_c_4_p N_VDD_c_71_n 0.0016649f
cc_5 N_VSS_c_5_p N_VDD_c_71_n 0.00583639f
cc_6 N_VSS_c_6_p N_VDD_c_71_n 0.00213268f
cc_7 N_VSS_c_7_p N_VDD_c_75_n 9.61646e-19
cc_8 N_VSS_c_8_p N_VDD_c_75_n 4.3619e-19
cc_9 N_VSS_c_5_p N_VDD_c_75_n 0.00351219f
cc_10 N_VSS_c_10_p N_VDD_c_75_n 0.00128683f
cc_11 N_VSS_c_4_p N_VDD_c_79_n 0.00221042f
cc_12 N_VSS_c_4_p N_VDD_c_80_n 7.48389e-19
cc_13 N_VSS_c_13_p N_VDD_c_81_n 0.00144388f
cc_14 N_VSS_c_14_p N_VDD_c_81_n 2.81922e-19
cc_15 N_VSS_c_7_p N_VDD_c_81_n 0.00161703f
cc_16 N_VSS_c_8_p N_VDD_c_81_n 2.03837e-19
cc_17 N_VSS_c_17_p N_VDD_c_81_n 0.00338232f
cc_18 N_VSS_c_18_p N_VDD_c_81_n 0.00635521f
cc_19 N_VSS_c_19_p N_VDD_c_81_n 7.61747e-19
cc_20 N_VSS_XI9.X0_PGS N_VDD_c_88_n 2.28184e-19
cc_21 N_VSS_XI2.X0_PGS N_VDD_c_88_n 2.56778e-19
cc_22 N_VSS_c_7_p N_VDD_c_88_n 5.65664e-19
cc_23 N_VSS_c_23_p N_VDD_c_88_n 0.00181281f
cc_24 N_VSS_c_8_p N_VDD_c_88_n 2.30125e-19
cc_25 N_VSS_c_25_p N_VDD_c_88_n 9.55109e-19
cc_26 N_VSS_c_2_p N_VDD_c_94_n 4.8598e-19
cc_27 N_VSS_c_23_p N_VDD_c_94_n 0.00161703f
cc_28 N_VSS_c_25_p N_VDD_c_94_n 2.03837e-19
cc_29 N_VSS_c_18_p N_VDD_c_94_n 0.00145178f
cc_30 N_VSS_c_30_p N_VDD_c_94_n 0.00590089f
cc_31 N_VSS_c_31_p N_VDD_c_94_n 7.74609e-19
cc_32 N_VSS_c_23_p N_VDD_c_100_n 8.94411e-19
cc_33 N_VSS_c_33_p N_VDD_c_100_n 3.85245e-19
cc_34 N_VSS_c_5_p N_VDD_c_102_n 0.00104993f
cc_35 N_VSS_c_18_p N_VDD_c_103_n 0.00119068f
cc_36 N_VSS_c_23_p N_VDD_c_104_n 3.48267e-19
cc_37 N_VSS_c_25_p N_VDD_c_104_n 8.0279e-19
cc_38 N_VSS_c_8_p N_A_c_156_n 0.00234241f
cc_39 N_VSS_c_7_p N_A_c_157_n 8.12473e-19
cc_40 N_VSS_c_8_p N_A_c_157_n 5.42695e-19
cc_41 N_VSS_c_5_p N_A_c_157_n 6.55807e-19
cc_42 N_VSS_c_42_p N_A_c_160_n 7.84334e-19
cc_43 N_VSS_c_7_p N_A_c_160_n 4.56568e-19
cc_44 N_VSS_c_8_p N_A_c_160_n 0.00184767f
cc_45 N_VSS_XI7.X0_S N_NET1_XI7.X0_D 3.43419e-19
cc_46 N_VSS_c_4_p N_NET1_XI7.X0_D 3.48267e-19
cc_47 N_VSS_c_25_p N_NET1_c_183_n 0.00413078f
cc_48 N_VSS_XI2.X0_PGD N_NET1_c_184_n 4.20799e-19
cc_49 N_VSS_c_49_p N_NET1_c_185_n 9.28737e-19
cc_50 N_VSS_c_25_p N_NET1_c_185_n 2.03369e-19
cc_51 N_VSS_XI7.X0_S N_NET1_c_187_n 3.48267e-19
cc_52 N_VSS_c_4_p N_NET1_c_187_n 8.46599e-19
cc_53 N_VSS_c_5_p N_NET1_c_187_n 2.07501e-19
cc_54 N_VSS_c_23_p N_NET1_c_190_n 0.00125323f
cc_55 N_VSS_c_25_p N_NET1_c_190_n 4.64764e-19
cc_56 N_VSS_c_5_p N_NET1_c_190_n 3.39684e-19
cc_57 N_VSS_c_23_p N_NET1_c_193_n 4.56568e-19
cc_58 N_VSS_c_25_p N_NET1_c_193_n 6.1245e-19
cc_59 N_VSS_c_5_p N_NET1_c_195_n 2.06399e-19
cc_60 N_VSS_c_18_p N_NET1_c_195_n 0.00149275f
cc_61 N_VSS_XI8.X0_PGD N_B_c_232_n 6.72196e-19
cc_62 N_VSS_XI9.X0_PGD N_B_c_232_n 6.72196e-19
cc_63 N_VSS_XI8.X0_PGS N_B_c_234_n 7.85613e-19
cc_64 N_VSS_XI1.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_65 N_VSS_c_65_p N_Z_XI2.X0_D 3.48267e-19
cc_66 N_VSS_c_65_p N_Z_c_260_n 5.37696e-19
cc_67 N_VSS_c_30_p N_Z_c_260_n 2.64173e-19
cc_68 N_VSS_c_68_p N_Z_c_260_n 2.7826e-19
cc_69 N_VDD_XI7.X0_PGD N_A_XI7.X0_CG 4.88425e-19
cc_70 N_VDD_c_79_n N_A_c_164_n 3.72495e-19
cc_71 N_VDD_c_71_n N_A_c_157_n 0.00273528f
cc_72 N_VDD_c_79_n N_A_c_157_n 7.03725e-19
cc_73 N_VDD_XI7.X0_PGD N_A_c_167_n 2.88617e-19
cc_74 N_VDD_c_71_n N_A_c_167_n 3.68786e-19
cc_75 N_VDD_c_79_n N_A_c_167_n 4.3265e-19
cc_76 N_VDD_c_113_p N_A_c_167_n 7.96439e-19
cc_77 N_VDD_c_71_n N_A_c_160_n 5.09899e-19
cc_78 N_VDD_c_79_n N_NET1_XI7.X0_D 9.18655e-19
cc_79 N_VDD_c_116_p N_NET1_XI7.X0_D 8.835e-19
cc_80 N_VDD_c_113_p N_NET1_XI7.X0_D 0.00132057f
cc_81 N_VDD_XI8.X0_S N_NET1_XI8.X0_D 3.43419e-19
cc_82 N_VDD_XI9.X0_S N_NET1_XI8.X0_D 3.43419e-19
cc_83 N_VDD_c_80_n N_NET1_XI8.X0_D 3.74351e-19
cc_84 N_VDD_c_81_n N_NET1_XI8.X0_D 3.7884e-19
cc_85 N_VDD_c_88_n N_NET1_XI8.X0_D 3.48267e-19
cc_86 N_VDD_c_104_n N_NET1_XI1.X0_CG 8.03148e-19
cc_87 N_VDD_XI1.X0_PGD N_NET1_c_184_n 4.25379e-19
cc_88 N_VDD_XI7.X0_PGD N_NET1_c_187_n 2.94751e-19
cc_89 N_VDD_XI8.X0_S N_NET1_c_187_n 3.48267e-19
cc_90 N_VDD_XI9.X0_S N_NET1_c_187_n 3.48267e-19
cc_91 N_VDD_c_128_p N_NET1_c_187_n 5.10453e-19
cc_92 N_VDD_c_71_n N_NET1_c_187_n 6.49505e-19
cc_93 N_VDD_c_79_n N_NET1_c_187_n 0.00151981f
cc_94 N_VDD_c_80_n N_NET1_c_187_n 8.1398e-19
cc_95 N_VDD_c_81_n N_NET1_c_187_n 5.36364e-19
cc_96 N_VDD_c_116_p N_NET1_c_187_n 0.00366419f
cc_97 N_VDD_c_88_n N_NET1_c_187_n 7.99681e-19
cc_98 N_VDD_c_113_p N_NET1_c_187_n 8.835e-19
cc_99 N_VDD_c_79_n N_NET1_c_195_n 3.89533e-19
cc_100 N_VDD_c_81_n N_NET1_c_195_n 3.69547e-19
cc_101 N_VDD_c_116_p N_NET1_c_195_n 4.83374e-19
cc_102 N_VDD_c_88_n N_NET1_c_195_n 4.34102e-19
cc_103 N_VDD_XI7.X0_PGD N_B_XI7.X0_PGS 0.00320719f
cc_104 N_VDD_c_71_n N_B_XI7.X0_PGS 6.17633e-19
cc_105 N_VDD_c_79_n N_B_XI7.X0_PGS 2.2956e-19
cc_106 N_VDD_c_143_p N_B_c_232_n 0.00973324f
cc_107 N_VDD_c_81_n N_B_c_239_n 4.48125e-19
cc_108 N_VDD_c_116_p N_B_c_239_n 4.13122e-19
cc_109 N_VDD_c_113_p N_B_c_239_n 0.00150022f
cc_110 N_VDD_c_81_n N_B_c_242_n 2.66883e-19
cc_111 N_VDD_c_116_p N_B_c_242_n 3.55986e-19
cc_112 N_VDD_c_113_p N_B_c_242_n 3.81676e-19
cc_113 N_VDD_XI9.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_114 N_VDD_c_88_n N_Z_XI2.X0_D 3.48267e-19
cc_115 N_VDD_c_94_n N_Z_XI2.X0_D 3.7884e-19
cc_116 N_VDD_XI9.X0_S N_Z_c_260_n 3.48267e-19
cc_117 N_VDD_c_88_n N_Z_c_260_n 7.06424e-19
cc_118 N_VDD_c_94_n N_Z_c_260_n 5.12447e-19
cc_119 N_A_c_157_n N_NET1_c_187_n 0.00751692f
cc_120 N_A_c_167_n N_NET1_c_187_n 9.57699e-19
cc_121 N_A_c_160_n N_NET1_c_187_n 9.18163e-19
cc_122 N_A_XI7.X0_CG N_B_XI7.X0_PGS 4.5346e-19
cc_123 N_A_c_167_n N_B_XI7.X0_PGS 5.70584e-19
cc_124 N_A_c_157_n N_B_c_232_n 2.1473e-19
cc_125 N_A_c_167_n N_B_c_232_n 0.0014179f
cc_126 N_A_c_160_n N_B_c_232_n 0.00112482f
cc_127 N_A_c_160_n N_B_c_239_n 9.27569e-19
cc_128 N_NET1_c_187_n N_B_c_232_n 7.63501e-19
cc_129 N_NET1_c_187_n N_B_c_239_n 9.91045e-19
cc_130 N_NET1_c_190_n N_B_c_239_n 3.63713e-19
cc_131 N_NET1_c_193_n N_B_c_239_n 0.00197331f
cc_132 N_NET1_c_187_n N_B_c_242_n 0.00142922f
cc_133 N_NET1_c_190_n N_B_c_242_n 3.90886e-19
cc_134 N_NET1_c_193_n N_B_c_242_n 3.48267e-19
*
.ends
*
*
.subckt AND2_HPNW1 A B Y VDD VSS
xgate (VSS VDD A B Y) G3_AND2_N1
.ends
*
* File: G2_AOI21_N1.pex.netlist
* Created: Mon Apr 11 11:24:15 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_AOI21_N1_VSS 2 4 6 8 19 25 38 43 48 57 66 67 69 77 78 79 83 84 86
+ 88 89 Vss
c53 89 Vss 4.28045e-19
c54 86 Vss 0.00420179f
c55 84 Vss 0.00142701f
c56 83 Vss 8.42815e-19
c57 79 Vss 0.00125695f
c58 78 Vss 4.66086e-19
c59 77 Vss 0.00243143f
c60 69 Vss 0.00100335f
c61 68 Vss 0.00135524f
c62 67 Vss 0.00884313f
c63 66 Vss 0.00244299f
c64 57 Vss 0.00663377f
c65 48 Vss 1.70165e-19
c66 43 Vss 0.00203396f
c67 38 Vss 0.00129403f
c68 25 Vss 0.0827803f
c69 19 Vss 0.034042f
c70 18 Vss 0.0688517f
c71 8 Vss 0.0810091f
c72 6 Vss 0.00226958f
c73 4 Vss 0.0797379f
c74 2 Vss 0.00290534f
r75 85 89 0.551426
r76 85 86 13.3371
r77 84 89 0.551426
r78 83 88 0.326149
r79 83 84 4.12618
r80 79 89 0.0828784
r81 77 86 0.652036
r82 77 78 4.33457
r83 73 78 0.652036
r84 67 88 0.326149
r85 67 68 15.1308
r86 66 69 0.655813
r87 65 68 0.652298
r88 65 66 4.12618
r89 48 79 1.82344
r90 43 57 1.16709
r91 43 73 2.16729
r92 38 69 1.82344
r93 25 57 0.238214
r94 23 25 2.04225
r95 20 23 0.0685365
r96 18 23 0.5835
r97 18 19 2.8008
r98 15 19 0.652036
r99 8 20 2.5674
r100 6 48 1.16709
r101 4 15 2.5674
r102 2 38 1.16709
.ends

.subckt PM_G2_AOI21_N1_VDD 2 4 6 8 10 45 46 48 50 54 56 57 58 63 65 67 68 74 Vss
c60 74 Vss 0.00498639f
c61 68 Vss 3.56526e-19
c62 65 Vss 0.00188744f
c63 63 Vss 0.00658029f
c64 58 Vss 0.00166035f
c65 57 Vss 6.17427e-19
c66 56 Vss 0.0030725f
c67 54 Vss 0.0015334f
c68 50 Vss 0.0128179f
c69 48 Vss 0.00148319f
c70 46 Vss 0.00118366f
c71 45 Vss 0.00509044f
c72 33 Vss 0.0307391f
c73 26 Vss 0.10055f
c74 22 Vss 0.0348457f
c75 21 Vss 0.0712517f
c76 10 Vss 0.00241752f
c77 8 Vss 0.0830779f
c78 6 Vss 0.0830019f
c79 4 Vss 0.00285737f
c80 2 Vss 0.0825892f
r81 64 68 0.551426
r82 64 65 4.16786
r83 63 68 0.551426
r84 62 63 13.2955
r85 58 68 0.0828784
r86 58 60 1.82344
r87 56 62 0.652298
r88 56 57 4.22534
r89 54 74 1.16709
r90 52 57 0.652298
r91 52 54 2.12561
r92 51 67 0.326018
r93 50 65 0.652036
r94 50 51 15.6711
r95 46 48 1.82344
r96 45 67 0.326018
r97 44 46 0.655813
r98 44 45 4.16786
r99 29 74 0.238214
r100 27 33 0.494161
r101 27 29 1.45875
r102 26 30 0.652036
r103 26 29 1.45875
r104 23 33 0.128424
r105 21 33 0.494161
r106 21 22 2.8008
r107 18 22 0.652036
r108 10 60 1.16709
r109 8 30 2.5674
r110 6 23 2.5674
r111 4 48 1.16709
r112 2 18 2.5674
.ends

.subckt PM_G2_AOI21_N1_B 2 4 20 23 29 Vss
c19 29 Vss 0.00607059f
c20 23 Vss 9.01834e-19
c21 20 Vss 0.0916059f
c22 16 Vss 0.0586024f
c23 4 Vss 0.0980254f
c24 2 Vss 0.320472f
r25 26 29 1.16709
r26 23 26 0.0833571
r27 18 20 2.04225
r28 16 29 0.197068
r29 13 16 1.2837
r30 10 20 0.0685365
r31 8 18 0.0685365
r32 7 13 0.0685365
r33 4 10 3.0342
r34 2 8 8.6358
r35 2 7 2.5674
.ends

.subckt PM_G2_AOI21_N1_C 2 4 6 17 24 28 31 35 38 42 45 58 Vss
c45 58 Vss 0.00118496f
c46 45 Vss 0.00482667f
c47 38 Vss 0.00276154f
c48 31 Vss 0.00515878f
c49 28 Vss 0.0945059f
c50 24 Vss 0.0559062f
c51 17 Vss 1.54762e-19
c52 6 Vss 0.178585f
c53 4 Vss 0.147123f
c54 2 Vss 0.0809403f
r55 54 58 0.652036
r56 38 58 5.16814
r57 38 42 0.0416786
r58 31 45 1.16709
r59 31 54 8.58579
r60 31 35 0.0416786
r61 26 28 2.04225
r62 24 45 0.197068
r63 21 24 1.2837
r64 18 28 0.0685365
r65 17 38 1.16709
r66 13 26 0.0685365
r67 13 17 2.8008
r68 10 21 0.0685365
r69 6 18 5.835
r70 4 17 3.0342
r71 2 10 2.5674
.ends

.subckt PM_G2_AOI21_N1_Z 2 4 30 33 Vss
c30 30 Vss 0.00225284f
c31 4 Vss 0.00143442f
c32 2 Vss 0.00153036f
r33 33 35 3.83443
r34 30 33 5.33486
r35 4 35 1.16709
r36 2 30 1.16709
.ends

.subckt PM_G2_AOI21_N1_A 2 4 10 11 13 14 15 20 24 28 31 Vss
c37 31 Vss 4.87906e-19
c38 28 Vss 4.59888e-19
c39 24 Vss 1.50097e-19
c40 20 Vss 0.0822806f
c41 18 Vss 0.0247918f
c42 15 Vss 0.032139f
c43 14 Vss 0.0725371f
c44 13 Vss 0.0312529f
c45 11 Vss 0.0345237f
c46 10 Vss 0.122163f
c47 2 Vss 0.188674f
r48 28 31 1.16709
r49 24 31 0.262036
r50 20 31 0.238214
r51 18 24 0.326018
r52 18 20 0.64185
r53 15 24 2.50905
r54 14 24 0.326018
r55 14 24 0.1167
r56 13 15 0.652036
r57 12 13 1.22535
r58 10 12 0.652036
r59 10 11 3.09255
r60 7 11 0.652036
r61 4 20 2.4507
r62 2 7 6.1851
.ends

.subckt G2_AOI21_N1  VSS VDD B C Z A
*
* A	A
* Z	Z
* C	C
* B	B
* VDD	VDD
* VSS	VSS
XI1.X0 N_Z_XI1.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_B_XI1.X0_PGS N_VSS_XI1.X0_S
+ TIGFET_HPNW1
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_C_XI6.X0_PGS N_VDD_XI6.X0_S
+ TIGFET_HPNW1
XI5.X0 N_Z_XI1.X0_D N_VDD_XI5.X0_PGD N_C_XI5.X0_CG N_VDD_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW1
XI7.X0 N_Z_XI6.X0_D N_VSS_XI7.X0_PGD N_A_XI7.X0_CG N_C_XI7.X0_PGS N_VDD_XI7.X0_S
+ TIGFET_HPNW1
*
x_PM_G2_AOI21_N1_VSS N_VSS_XI1.X0_S N_VSS_XI6.X0_PGD N_VSS_XI5.X0_S
+ N_VSS_XI7.X0_PGD N_VSS_c_3_p N_VSS_c_46_p N_VSS_c_2_p N_VSS_c_4_p N_VSS_c_8_p
+ N_VSS_c_20_p N_VSS_c_23_p N_VSS_c_9_p N_VSS_c_1_p N_VSS_c_5_p N_VSS_c_6_p
+ N_VSS_c_13_p N_VSS_c_10_p N_VSS_c_16_p N_VSS_c_17_p VSS N_VSS_c_18_p Vss
+ PM_G2_AOI21_N1_VSS
x_PM_G2_AOI21_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI6.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI5.X0_PGS N_VDD_XI7.X0_S N_VDD_c_89_p N_VDD_c_54_n N_VDD_c_55_n
+ N_VDD_c_56_n N_VDD_c_77_p N_VDD_c_60_n N_VDD_c_64_n N_VDD_c_65_n N_VDD_c_67_n
+ N_VDD_c_72_n VDD N_VDD_c_75_n N_VDD_c_78_p Vss PM_G2_AOI21_N1_VDD
x_PM_G2_AOI21_N1_B N_B_XI1.X0_PGS N_B_XI6.X0_CG N_B_c_122_p B N_B_c_119_n Vss
+ PM_G2_AOI21_N1_B
x_PM_G2_AOI21_N1_C N_C_XI6.X0_PGS N_C_XI5.X0_CG N_C_XI7.X0_PGS N_C_c_143_n
+ N_C_c_146_n N_C_c_147_n N_C_c_134_n C N_C_c_136_n C N_C_c_137_n N_C_c_140_n
+ Vss PM_G2_AOI21_N1_C
x_PM_G2_AOI21_N1_Z N_Z_XI1.X0_D N_Z_XI6.X0_D N_Z_c_182_n Z Vss PM_G2_AOI21_N1_Z
x_PM_G2_AOI21_N1_A N_A_XI1.X0_CG N_A_XI7.X0_CG N_A_c_208_n N_A_c_225_n
+ N_A_c_226_n N_A_c_209_n N_A_c_227_n N_A_c_211_n N_A_c_212_n A N_A_c_216_n Vss
+ PM_G2_AOI21_N1_A
cc_1 N_VSS_c_1_p N_VDD_c_54_n 4.93612e-19
cc_2 N_VSS_c_2_p N_VDD_c_55_n 9.30121e-19
cc_3 N_VSS_c_3_p N_VDD_c_56_n 0.0011834f
cc_4 N_VSS_c_4_p N_VDD_c_56_n 0.00161703f
cc_5 N_VSS_c_5_p N_VDD_c_56_n 0.00445263f
cc_6 N_VSS_c_6_p N_VDD_c_56_n 0.00169823f
cc_7 N_VSS_XI5.X0_S N_VDD_c_60_n 3.83684e-19
cc_8 N_VSS_c_8_p N_VDD_c_60_n 4.79306e-19
cc_9 N_VSS_c_9_p N_VDD_c_60_n 0.0035571f
cc_10 N_VSS_c_10_p N_VDD_c_60_n 0.00109026f
cc_11 N_VSS_c_9_p N_VDD_c_64_n 0.00162315f
cc_12 N_VSS_c_8_p N_VDD_c_65_n 2.13058e-19
cc_13 N_VSS_c_13_p N_VDD_c_65_n 5.33968e-19
cc_14 N_VSS_XI5.X0_S N_VDD_c_67_n 9.5668e-19
cc_15 N_VSS_c_8_p N_VDD_c_67_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_67_n 0.00300233f
cc_17 N_VSS_c_17_p N_VDD_c_67_n 0.00605714f
cc_18 N_VSS_c_18_p N_VDD_c_67_n 8.91588e-19
cc_19 N_VSS_c_4_p N_VDD_c_72_n 4.42697e-19
cc_20 N_VSS_c_20_p N_VDD_c_72_n 3.70842e-19
cc_21 N_VSS_c_17_p N_VDD_c_72_n 0.00278561f
cc_22 N_VSS_c_17_p N_VDD_c_75_n 9.45256e-19
cc_23 N_VSS_c_23_p B 3.22996e-19
cc_24 N_VSS_c_9_p B 3.31649e-19
cc_25 N_VSS_XI6.X0_PGD N_C_XI6.X0_PGS 0.00161425f
cc_26 N_VSS_c_4_p N_C_c_134_n 5.88052e-19
cc_27 N_VSS_c_17_p N_C_c_134_n 0.00138265f
cc_28 N_VSS_c_17_p N_C_c_136_n 3.65158e-19
cc_29 N_VSS_XI6.X0_PGD N_C_c_137_n 3.23173e-19
cc_30 N_VSS_c_4_p N_C_c_137_n 3.44698e-19
cc_31 N_VSS_c_20_p N_C_c_137_n 3.34921e-19
cc_32 N_VSS_c_9_p N_C_c_140_n 0.00303126f
cc_33 N_VSS_c_17_p N_C_c_140_n 3.90377e-19
cc_34 N_VSS_XI1.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_35 N_VSS_XI5.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_XI1.X0_D 3.48267e-19
cc_37 N_VSS_c_8_p N_Z_XI1.X0_D 3.48267e-19
cc_38 N_VSS_XI1.X0_S N_Z_c_182_n 3.48267e-19
cc_39 N_VSS_XI5.X0_S N_Z_c_182_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_182_n 5.69026e-19
cc_41 N_VSS_c_8_p N_Z_c_182_n 5.69026e-19
cc_42 N_VSS_c_9_p N_Z_c_182_n 4.18012e-19
cc_43 N_VSS_c_17_p N_Z_c_182_n 5.20852e-19
cc_44 N_VSS_XI6.X0_PGD N_A_c_208_n 7.38139e-19
cc_45 N_VSS_XI7.X0_PGD N_A_c_209_n 0.00160007f
cc_46 N_VSS_c_46_p N_A_c_209_n 3.07681e-19
cc_47 N_VSS_c_20_p N_A_c_211_n 0.00255152f
cc_48 N_VSS_c_46_p N_A_c_212_n 8.89952e-19
cc_49 N_VSS_c_20_p N_A_c_212_n 2.75949e-19
cc_50 N_VSS_c_4_p A 5.37794e-19
cc_51 N_VSS_c_20_p A 4.56568e-19
cc_52 N_VSS_c_4_p N_A_c_216_n 4.56568e-19
cc_53 N_VSS_c_20_p N_A_c_216_n 6.1245e-19
cc_54 N_VDD_XI1.X0_PGD N_B_XI1.X0_PGS 0.0015605f
cc_55 N_VDD_c_77_p B 5.21626e-19
cc_56 N_VDD_c_78_p B 3.48267e-19
cc_57 N_VDD_XI1.X0_PGD N_B_c_119_n 3.73456e-19
cc_58 N_VDD_c_77_p N_B_c_119_n 4.2695e-19
cc_59 N_VDD_c_78_p N_B_c_119_n 5.71625e-19
cc_60 N_VDD_c_78_p N_C_XI5.X0_CG 0.00117555f
cc_61 N_VDD_c_77_p N_C_c_143_n 4.85469e-19
cc_62 N_VDD_c_67_n N_C_c_143_n 5.82627e-19
cc_63 N_VDD_c_78_p N_C_c_143_n 0.00182135f
cc_64 N_VDD_c_56_n N_C_c_146_n 3.54083e-19
cc_65 N_VDD_XI5.X0_PGS N_C_c_147_n 7.91098e-19
cc_66 N_VDD_c_67_n N_C_c_147_n 4.33233e-19
cc_67 N_VDD_c_89_p N_C_c_134_n 3.48763e-19
cc_68 N_VDD_c_55_n N_C_c_134_n 3.25844e-19
cc_69 N_VDD_c_56_n N_C_c_134_n 0.00156477f
cc_70 N_VDD_c_56_n N_C_c_136_n 7.40864e-19
cc_71 N_VDD_c_77_p N_C_c_136_n 5.82566e-19
cc_72 N_VDD_c_67_n N_C_c_136_n 4.90875e-19
cc_73 N_VDD_c_78_p N_C_c_136_n 4.56568e-19
cc_74 N_VDD_c_89_p N_C_c_137_n 4.55865e-19
cc_75 N_VDD_c_56_n N_C_c_137_n 2.55177e-19
cc_76 N_VDD_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_77 N_VDD_XI7.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_78 N_VDD_c_55_n N_Z_XI6.X0_D 3.72199e-19
cc_79 N_VDD_c_56_n N_Z_XI6.X0_D 3.7884e-19
cc_80 N_VDD_c_65_n N_Z_XI6.X0_D 3.72199e-19
cc_81 N_VDD_XI6.X0_S N_Z_c_182_n 3.48267e-19
cc_82 N_VDD_XI7.X0_S N_Z_c_182_n 3.48267e-19
cc_83 N_VDD_c_55_n N_Z_c_182_n 5.68773e-19
cc_84 N_VDD_c_56_n N_Z_c_182_n 6.9352e-19
cc_85 N_VDD_c_65_n N_Z_c_182_n 7.77875e-19
cc_86 N_VDD_c_67_n N_Z_c_182_n 9.95668e-19
cc_87 N_VDD_XI1.X0_PGD N_A_c_208_n 6.1925e-19
cc_88 N_VDD_XI5.X0_PGD N_A_c_209_n 3.67852e-19
cc_89 N_VDD_c_67_n A 3.35548e-19
cc_90 N_VDD_c_56_n N_A_c_216_n 2.29043e-19
cc_91 N_VDD_c_67_n N_A_c_216_n 3.66936e-19
cc_92 N_B_c_122_p N_C_XI6.X0_PGS 0.00189436f
cc_93 N_B_XI1.X0_PGS N_C_XI5.X0_CG 2.46172e-19
cc_94 N_B_c_122_p N_C_XI7.X0_PGS 4.95875e-19
cc_95 N_B_c_122_p N_C_c_146_n 3.12087e-19
cc_96 N_B_XI1.X0_PGS N_Z_c_182_n 2.61881e-19
cc_97 N_B_XI1.X0_PGS N_A_XI1.X0_CG 0.00900711f
cc_98 N_B_c_119_n N_A_XI1.X0_CG 0.00150571f
cc_99 N_B_c_122_p N_A_c_225_n 0.00163406f
cc_100 N_B_XI1.X0_PGS N_A_c_226_n 6.07734e-19
cc_101 N_B_c_122_p N_A_c_227_n 0.00136506f
cc_102 N_B_c_122_p N_A_c_216_n 2.87722e-19
cc_103 N_C_c_143_n N_Z_c_182_n 9.29334e-19
cc_104 N_C_c_134_n N_Z_c_182_n 0.00223036f
cc_105 N_C_c_136_n N_Z_c_182_n 0.00299789f
cc_106 N_C_c_140_n N_Z_c_182_n 2.70867e-19
cc_107 N_C_XI5.X0_CG N_A_XI1.X0_CG 5.49495e-19
cc_108 N_C_c_143_n N_A_XI1.X0_CG 5.65259e-19
cc_109 N_C_XI7.X0_PGS N_A_c_208_n 8.10159e-19
cc_110 N_C_c_147_n N_A_c_208_n 0.00121323f
cc_111 N_C_XI7.X0_PGS N_A_c_211_n 5.00154e-19
cc_112 N_C_c_143_n N_A_c_212_n 9.55393e-19
cc_113 N_C_c_143_n A 4.56568e-19
cc_114 N_C_c_136_n A 6.2998e-19
cc_115 N_C_XI7.X0_PGS N_A_c_216_n 0.00570455f
cc_116 N_C_c_143_n N_A_c_216_n 8.77002e-19
cc_117 N_C_c_147_n N_A_c_216_n 0.00119367f
cc_118 N_C_c_136_n N_A_c_216_n 4.56568e-19
cc_119 N_Z_c_182_n N_A_XI1.X0_CG 5.75111e-19
cc_120 N_Z_c_182_n N_A_c_208_n 4.34888e-19
cc_121 N_Z_c_182_n A 0.0015179f
cc_122 N_Z_c_182_n N_A_c_216_n 8.99071e-19
*
.ends
*
*
.subckt AOI21_HPNW1 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 B0 Y A0) G2_AOI21_N1
.ends
*
* File: G2_BUF1_N1.pex.netlist
* Created: Wed Mar  2 15:26:00 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_BUF1_N1_VDD 2 4 7 11 28 32 52 56 58 59 63 67 69 73 77 90 95 Vss
c58 95 Vss 0.00471589f
c59 90 Vss 0.0048335f
c60 80 Vss 7.0893e-19
c61 79 Vss 7.0893e-19
c62 77 Vss 0.00107913f
c63 73 Vss 0.00106523f
c64 70 Vss 0.00175834f
c65 69 Vss 0.00726612f
c66 67 Vss 0.00110053f
c67 63 Vss 0.00110053f
c68 60 Vss 0.00175834f
c69 59 Vss 0.00712138f
c70 58 Vss 0.00330526f
c71 56 Vss 0.00424287f
c72 52 Vss 0.00330526f
c73 32 Vss 0.0346129f
c74 31 Vss 0.101192f
c75 28 Vss 0.0346129f
c76 27 Vss 0.101192f
c77 11 Vss 0.16682f
c78 7 Vss 0.16682f
c79 4 Vss 0.00203161f
c80 2 Vss 0.00233151f
r81 77 95 1.16709
r82 75 77 2.16729
r83 73 90 1.16709
r84 71 73 2.16729
r85 69 75 0.652036
r86 69 70 10.1279
r87 65 80 0.0828784
r88 65 67 1.82344
r89 61 79 0.0828784
r90 61 63 1.82344
r91 59 71 0.652036
r92 59 60 10.1279
r93 58 70 0.652036
r94 57 80 0.551426
r95 57 58 4.16786
r96 54 80 0.551426
r97 54 56 3.45932
r98 53 79 0.551426
r99 53 56 1.45875
r100 52 79 0.551426
r101 51 60 0.652036
r102 51 52 4.16786
r103 34 95 0.238214
r104 32 34 1.45875
r105 31 38 0.652036
r106 31 34 1.45875
r107 30 90 0.238214
r108 28 30 1.45875
r109 27 35 0.652036
r110 27 30 1.45875
r111 24 32 0.652036
r112 21 28 0.652036
r113 11 38 2.5674
r114 11 24 2.5674
r115 7 35 2.5674
r116 7 21 2.5674
r117 4 67 1.16709
r118 2 63 1.16709
.ends

.subckt PM_G2_BUF1_N1_VSS 3 7 10 12 27 28 31 32 52 57 62 67 72 77 97 98 99 100
+ 101 105 110 114 116 Vss
c60 118 Vss 6.78504e-19
c61 117 Vss 6.78504e-19
c62 116 Vss 0.00235663f
c63 114 Vss 0.00287691f
c64 110 Vss 0.00235663f
c65 105 Vss 9.66804e-19
c66 101 Vss 8.0746e-19
c67 100 Vss 5.83649e-19
c68 99 Vss 0.00631424f
c69 98 Vss 5.83649e-19
c70 97 Vss 0.00625937f
c71 77 Vss 0.00398915f
c72 72 Vss 0.00399741f
c73 67 Vss 1.62164e-19
c74 62 Vss 3.56438e-22
c75 57 Vss 8.13664e-19
c76 52 Vss 7.92706e-19
c77 34 Vss 1.28632e-19
c78 32 Vss 0.0341976f
c79 31 Vss 0.0984533f
c80 28 Vss 0.0341976f
c81 27 Vss 0.0984533f
c82 12 Vss 0.00237948f
c83 10 Vss 0.00207958f
c84 7 Vss 0.16682f
c85 3 Vss 0.16682f
r86 115 118 0.551426
r87 115 116 4.16786
r88 112 118 0.551426
r89 112 114 2.12561
r90 111 117 0.551426
r91 111 114 2.79246
r92 110 117 0.551426
r93 109 110 4.16786
r94 105 118 0.0828784
r95 101 117 0.0828784
r96 99 116 0.652036
r97 99 100 10.1279
r98 97 109 0.652036
r99 97 98 10.1279
r100 93 100 0.652036
r101 89 98 0.652036
r102 67 105 1.82344
r103 62 101 1.82344
r104 57 77 1.16709
r105 57 93 2.16729
r106 52 72 1.16709
r107 52 89 2.16729
r108 34 77 0.238214
r109 32 34 1.45875
r110 31 38 0.652036
r111 31 34 1.45875
r112 30 72 0.238214
r113 28 30 1.45875
r114 27 35 0.652036
r115 27 30 1.45875
r116 24 32 0.652036
r117 21 28 0.652036
r118 12 67 1.16709
r119 10 62 1.16709
r120 7 38 2.5674
r121 7 24 2.5674
r122 3 35 2.5674
r123 3 21 2.5674
.ends

.subckt PM_G2_BUF1_N1_A 2 4 9 12 22 25 28 Vss
c18 28 Vss 0.00276471f
c19 25 Vss 3.55586e-19
c20 12 Vss 0.20721f
c21 9 Vss 0.0715834f
c22 7 Vss 0.0247918f
c23 4 Vss 0.0847975f
r24 25 28 1.16709
r25 22 25 0.0795682
r26 15 28 0.0476429
r27 13 15 0.326018
r28 13 15 0.1167
r29 12 16 0.652036
r30 12 15 6.7686
r31 9 28 0.357321
r32 7 15 0.326018
r33 7 9 0.40845
r34 4 16 2.5674
r35 2 9 2.15895
.ends

.subckt PM_G2_BUF1_N1_Z 2 19 Vss
c15 19 Vss 2.80869e-19
c16 2 Vss 0.00176567f
r17 16 19 0.0364688
r18 2 16 1.16709
.ends

.subckt PM_G2_BUF1_N1_NET17 2 4 6 18 36 41 50 58 Vss
c37 58 Vss 5.85801e-19
c38 50 Vss 0.00307045f
c39 41 Vss 0.0013766f
c40 36 Vss 0.00137137f
c41 22 Vss 0.0247918f
c42 19 Vss 0.0295882f
c43 18 Vss 0.176231f
c44 6 Vss 0.0715834f
c45 4 Vss 0.00176567f
c46 2 Vss 0.0847975f
r47 54 58 0.653045
r48 41 50 1.16709
r49 41 58 2.1395
r50 36 54 3.45932
r51 28 50 0.0476429
r52 26 50 0.357321
r53 22 28 0.326018
r54 22 26 0.40845
r55 19 28 6.7686
r56 18 28 0.326018
r57 18 28 0.1167
r58 15 19 0.652036
r59 6 26 2.15895
r60 4 36 1.16709
r61 2 15 2.5674
.ends

.subckt G2_BUF1_N1  VDD VSS A Z
*
* Z	Z
* A	A
* VSS	VSS
* VDD	VDD
XI3.X0 N_Z_XI3.X0_D N_VSS_XI3.X0_PGD N_NET17_XI3.X0_CG N_VSS_XI3.X0_PGD
+ N_VDD_XI3.X0_S TIGFET_HPNW1
XI2.X0 N_NET17_XI2.X0_D N_VSS_XI2.X0_PGD N_A_XI2.X0_CG N_VSS_XI2.X0_PGD
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI0.X0 N_Z_XI3.X0_D N_VDD_XI0.X0_PGD N_NET17_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW1
XI1.X0 N_NET17_XI2.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW1
*
x_PM_G2_BUF1_N1_VDD N_VDD_XI3.X0_S N_VDD_XI2.X0_S N_VDD_XI0.X0_PGD
+ N_VDD_XI1.X0_PGD N_VDD_c_3_p N_VDD_c_6_p N_VDD_c_9_p VDD N_VDD_c_13_p
+ N_VDD_c_4_p N_VDD_c_38_p N_VDD_c_43_p N_VDD_c_7_p N_VDD_c_11_p N_VDD_c_15_p
+ N_VDD_c_12_p N_VDD_c_16_p Vss PM_G2_BUF1_N1_VDD
x_PM_G2_BUF1_N1_VSS N_VSS_XI3.X0_PGD N_VSS_XI2.X0_PGD N_VSS_XI0.X0_S
+ N_VSS_XI1.X0_S N_VSS_c_61_n N_VSS_c_63_n N_VSS_c_64_n N_VSS_c_66_n
+ N_VSS_c_67_n N_VSS_c_71_n N_VSS_c_101_p N_VSS_c_110_p N_VSS_c_75_n
+ N_VSS_c_79_n N_VSS_c_83_n N_VSS_c_84_n N_VSS_c_85_n N_VSS_c_86_n N_VSS_c_104_p
+ N_VSS_c_112_p N_VSS_c_87_n VSS N_VSS_c_88_n Vss PM_G2_BUF1_N1_VSS
x_PM_G2_BUF1_N1_A N_A_XI2.X0_CG N_A_XI1.X0_CG N_A_c_124_n N_A_c_120_n A
+ N_A_c_122_n N_A_c_123_n Vss PM_G2_BUF1_N1_A
x_PM_G2_BUF1_N1_Z N_Z_XI3.X0_D Z Vss PM_G2_BUF1_N1_Z
x_PM_G2_BUF1_N1_NET17 N_NET17_XI3.X0_CG N_NET17_XI2.X0_D N_NET17_XI0.X0_CG
+ N_NET17_c_155_n N_NET17_c_157_n N_NET17_c_160_n N_NET17_c_164_n
+ N_NET17_c_168_n Vss PM_G2_BUF1_N1_NET17
cc_1 N_VDD_XI0.X0_PGD N_VSS_XI3.X0_PGD 0.00173038f
cc_2 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00173038f
cc_3 N_VDD_c_3_p N_VSS_c_61_n 0.00173038f
cc_4 N_VDD_c_4_p N_VSS_c_61_n 2.91357e-19
cc_5 N_VDD_c_4_p N_VSS_c_63_n 3.24852e-19
cc_6 N_VDD_c_6_p N_VSS_c_64_n 0.00173038f
cc_7 N_VDD_c_7_p N_VSS_c_64_n 2.91357e-19
cc_8 N_VDD_c_7_p N_VSS_c_66_n 3.24852e-19
cc_9 N_VDD_c_9_p N_VSS_c_67_n 8.69498e-19
cc_10 N_VDD_c_4_p N_VSS_c_67_n 0.00141228f
cc_11 N_VDD_c_11_p N_VSS_c_67_n 0.00106872f
cc_12 N_VDD_c_12_p N_VSS_c_67_n 3.48267e-19
cc_13 N_VDD_c_13_p N_VSS_c_71_n 8.69498e-19
cc_14 N_VDD_c_7_p N_VSS_c_71_n 0.00141228f
cc_15 N_VDD_c_15_p N_VSS_c_71_n 0.00106872f
cc_16 N_VDD_c_16_p N_VSS_c_71_n 3.48267e-19
cc_17 N_VDD_c_9_p N_VSS_c_75_n 3.66936e-19
cc_18 N_VDD_c_4_p N_VSS_c_75_n 0.00112249f
cc_19 N_VDD_c_11_p N_VSS_c_75_n 3.99794e-19
cc_20 N_VDD_c_12_p N_VSS_c_75_n 8.09245e-19
cc_21 N_VDD_c_13_p N_VSS_c_79_n 3.66936e-19
cc_22 N_VDD_c_7_p N_VSS_c_79_n 0.00112249f
cc_23 N_VDD_c_15_p N_VSS_c_79_n 3.99794e-19
cc_24 N_VDD_c_16_p N_VSS_c_79_n 8.09245e-19
cc_25 N_VDD_c_4_p N_VSS_c_83_n 0.00554293f
cc_26 N_VDD_c_4_p N_VSS_c_84_n 0.0017359f
cc_27 N_VDD_c_7_p N_VSS_c_85_n 0.00562924f
cc_28 N_VDD_c_7_p N_VSS_c_86_n 0.0017359f
cc_29 N_VDD_c_11_p N_VSS_c_87_n 3.85245e-19
cc_30 N_VDD_c_15_p N_VSS_c_88_n 3.85245e-19
cc_31 N_VDD_c_16_p N_A_XI1.X0_CG 0.00254294f
cc_32 N_VDD_XI0.X0_PGD N_A_c_120_n 4.08785e-19
cc_33 N_VDD_XI1.X0_PGD N_A_c_120_n 4.04053e-19
cc_34 VDD N_A_c_122_n 5.94555e-19
cc_35 VDD N_A_c_123_n 4.56718e-19
cc_36 N_VDD_XI3.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_37 N_VDD_c_4_p N_Z_XI3.X0_D 3.7884e-19
cc_38 N_VDD_c_38_p N_Z_XI3.X0_D 3.72199e-19
cc_39 N_VDD_XI3.X0_S Z 3.48267e-19
cc_40 N_VDD_c_4_p Z 5.12447e-19
cc_41 N_VDD_c_38_p Z 7.4527e-19
cc_42 N_VDD_XI2.X0_S N_NET17_XI2.X0_D 3.43419e-19
cc_43 N_VDD_c_43_p N_NET17_XI2.X0_D 3.72199e-19
cc_44 N_VDD_c_12_p N_NET17_XI0.X0_CG 0.0023817f
cc_45 N_VDD_XI0.X0_PGD N_NET17_c_155_n 4.04053e-19
cc_46 N_VDD_XI1.X0_PGD N_NET17_c_155_n 4.08785e-19
cc_47 N_VDD_XI2.X0_S N_NET17_c_157_n 3.48267e-19
cc_48 N_VDD_c_43_p N_NET17_c_157_n 8.0086e-19
cc_49 N_VDD_c_7_p N_NET17_c_157_n 5.01863e-19
cc_50 N_VDD_c_11_p N_NET17_c_160_n 6.85072e-19
cc_51 N_VDD_c_15_p N_NET17_c_160_n 3.98507e-19
cc_52 N_VDD_c_12_p N_NET17_c_160_n 4.99367e-19
cc_53 N_VDD_c_16_p N_NET17_c_160_n 3.0441e-19
cc_54 N_VDD_c_11_p N_NET17_c_164_n 4.85469e-19
cc_55 N_VDD_c_15_p N_NET17_c_164_n 3.00204e-19
cc_56 N_VDD_c_12_p N_NET17_c_164_n 0.0014909f
cc_57 N_VDD_c_16_p N_NET17_c_164_n 6.61247e-19
cc_58 VDD N_NET17_c_168_n 3.1911e-19
cc_59 N_VSS_c_79_n N_A_c_124_n 0.0023454f
cc_60 N_VSS_XI3.X0_PGD N_A_c_120_n 4.07282e-19
cc_61 N_VSS_XI2.X0_PGD N_A_c_120_n 3.99472e-19
cc_62 N_VSS_c_67_n N_A_c_122_n 2.85158e-19
cc_63 N_VSS_c_71_n N_A_c_122_n 5.53028e-19
cc_64 N_VSS_c_75_n N_A_c_122_n 3.0441e-19
cc_65 N_VSS_c_79_n N_A_c_122_n 4.99367e-19
cc_66 N_VSS_c_67_n N_A_c_123_n 2.82333e-19
cc_67 N_VSS_c_71_n N_A_c_123_n 4.56568e-19
cc_68 N_VSS_c_75_n N_A_c_123_n 6.61247e-19
cc_69 N_VSS_c_79_n N_A_c_123_n 0.0014909f
cc_70 N_VSS_XI0.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_71 N_VSS_c_101_p N_Z_XI3.X0_D 3.48267e-19
cc_72 N_VSS_XI0.X0_S Z 3.48267e-19
cc_73 N_VSS_c_101_p Z 4.99861e-19
cc_74 N_VSS_c_104_p Z 2.7826e-19
cc_75 N_VSS_c_75_n N_NET17_XI3.X0_CG 0.00250664f
cc_76 N_VSS_XI1.X0_S N_NET17_XI2.X0_D 3.43419e-19
cc_77 N_VSS_XI3.X0_PGD N_NET17_c_155_n 3.99472e-19
cc_78 N_VSS_XI2.X0_PGD N_NET17_c_155_n 4.07282e-19
cc_79 N_VSS_XI1.X0_S N_NET17_c_157_n 3.48267e-19
cc_80 N_VSS_c_110_p N_NET17_c_157_n 4.8288e-19
cc_81 N_VSS_c_85_n N_NET17_c_157_n 5.36354e-19
cc_82 N_VSS_c_112_p N_NET17_c_157_n 5.49885e-19
cc_83 VSS N_NET17_c_157_n 6.44069e-19
cc_84 N_VSS_c_83_n N_NET17_c_160_n 3.16821e-19
cc_85 N_VSS_c_85_n N_NET17_c_160_n 2.03753e-19
cc_86 VSS N_NET17_c_160_n 8.09756e-19
cc_87 N_VSS_c_83_n N_NET17_c_168_n 0.00101305f
cc_88 N_VSS_c_85_n N_NET17_c_168_n 5.70583e-19
cc_89 N_A_c_120_n N_NET17_c_155_n 0.00954069f
cc_90 N_A_c_122_n N_NET17_c_157_n 8.44937e-19
cc_91 N_Z_XI3.X0_D N_NET17_XI2.X0_D 2.56268e-19
cc_92 Z N_NET17_XI2.X0_D 3.17139e-19
cc_93 N_Z_XI3.X0_D N_NET17_c_157_n 3.17139e-19
cc_94 Z N_NET17_c_157_n 3.16516e-19
*
.ends
*
*
.subckt BUF1_HPNW1 A Y VDD VSS
xgate (VDD VSS A Y) G2_BUF1_N1
.ends
*
* File: G3_DFFQ1_N1.pex.netlist
* Created: Tue Apr  5 22:58:19 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_DFFQ1_N1_VSS 2 4 6 8 10 12 14 29 42 44 49 67 72 78 83 88 93 102
+ 111 116 125 126 127 128 132 137 142 148 154 156 161 163 165 166 167 Vss
c117 167 Vss 4.28045e-19
c118 166 Vss 3.75522e-19
c119 165 Vss 3.75522e-19
c120 164 Vss 6.13404e-19
c121 163 Vss 0.00437039f
c122 161 Vss 0.00140798f
c123 156 Vss 0.00134457f
c124 154 Vss 0.0025067f
c125 148 Vss 0.00439094f
c126 142 Vss 0.00297776f
c127 132 Vss 0.00193747f
c128 128 Vss 7.01403e-19
c129 127 Vss 8.12244e-19
c130 126 Vss 0.00567951f
c131 125 Vss 0.00148961f
c132 116 Vss 0.00596988f
c133 111 Vss 0.00418189f
c134 102 Vss 0.00407665f
c135 93 Vss 1.70165e-19
c136 88 Vss 0.00119073f
c137 83 Vss 5.15444e-19
c138 78 Vss 0.00173585f
c139 72 Vss 0.00866259f
c140 67 Vss 0.00134806f
c141 49 Vss 0.0560391f
c142 44 Vss 0.0560391f
c143 42 Vss 7.82991e-20
c144 29 Vss 0.0355813f
c145 28 Vss 0.101268f
c146 14 Vss 0.0832368f
c147 12 Vss 0.00370216f
c148 10 Vss 0.0027334f
c149 8 Vss 0.0822683f
c150 6 Vss 0.0792534f
c151 4 Vss 0.0793599f
c152 2 Vss 0.00198471f
r153 162 167 0.551426
r154 162 163 13.3371
r155 161 167 0.551426
r156 160 161 4.16786
r157 156 167 0.0828784
r158 155 166 0.494161
r159 154 163 0.652036
r160 154 155 4.37625
r161 150 166 0.128424
r162 149 165 0.494161
r163 148 160 0.652036
r164 148 149 10.1279
r165 144 165 0.128424
r166 143 164 0.494161
r167 142 166 0.494161
r168 142 143 7.46046
r169 138 164 0.128424
r170 132 164 0.494161
r171 132 137 1.00029
r172 126 165 0.494161
r173 126 127 15.8795
r174 125 128 0.655813
r175 124 127 0.652036
r176 124 125 4.16786
r177 93 156 1.82344
r178 88 116 1.16709
r179 88 150 2.16729
r180 83 111 1.16709
r181 83 144 2.16729
r182 78 138 4.83471
r183 75 137 1.29204
r184 72 102 1.16709
r185 72 75 12.4202
r186 67 128 1.82344
r187 49 116 0.197068
r188 46 49 1.2837
r189 42 111 0.197068
r190 42 44 1.2837
r191 38 46 0.0685365
r192 35 44 0.0685365
r193 31 102 0.0476429
r194 29 31 1.45875
r195 28 32 0.652036
r196 28 31 1.45875
r197 25 29 0.652036
r198 14 38 2.5674
r199 12 93 1.16709
r200 10 78 1.16709
r201 8 35 2.5674
r202 6 32 2.5674
r203 4 25 2.5674
r204 2 67 1.16709
.ends

.subckt PM_G3_DFFQ1_N1_CK 2 4 6 8 18 25 37 40 Vss
c31 40 Vss 0.00572916f
c32 37 Vss 3.65059e-19
c33 33 Vss 0.0299355f
c34 25 Vss 0.165118f
c35 18 Vss 0.186407f
c36 15 Vss 0.077884f
c37 13 Vss 0.0247918f
c38 6 Vss 0.441644f
c39 4 Vss 0.0840059f
r40 37 40 1.16709
r41 26 33 0.494161
r42 25 27 0.652036
r43 25 26 4.84305
r44 22 33 0.128424
r45 21 40 0.238214
r46 19 21 0.326018
r47 19 21 0.1167
r48 18 33 0.494161
r49 18 21 6.7686
r50 15 21 0.262036
r51 13 21 0.326018
r52 13 15 0.05835
r53 6 8 12.837
r54 6 27 2.5674
r55 4 22 2.5674
r56 2 15 2.50905
.ends

.subckt PM_G3_DFFQ1_N1_VDD 2 4 6 10 12 14 28 42 44 49 63 64 65 70 72 76 78 79 82
+ 84 86 91 93 95 96 98 99 100 102 104 113 118 Vss
c117 118 Vss 0.00660773f
c118 113 Vss 0.00546672f
c119 104 Vss 0.00477384f
c120 100 Vss 3.56526e-19
c121 99 Vss 2.39889e-19
c122 98 Vss 4.42156e-19
c123 96 Vss 0.00351049f
c124 95 Vss 5.22595e-19
c125 93 Vss 0.00279817f
c126 91 Vss 0.00684574f
c127 86 Vss 0.00166444f
c128 84 Vss 0.00296655f
c129 82 Vss 0.00146489f
c130 79 Vss 4.90412e-19
c131 78 Vss 0.00554983f
c132 76 Vss 5.91088e-19
c133 72 Vss 0.00336584f
c134 70 Vss 0.00240239f
c135 67 Vss 0.00178747f
c136 65 Vss 8.63831e-19
c137 64 Vss 0.00713032f
c138 63 Vss 0.00360153f
c139 49 Vss 0.0578141f
c140 44 Vss 0.0572437f
c141 42 Vss 7.44761e-20
c142 29 Vss 0.0373466f
c143 28 Vss 0.100964f
c144 14 Vss 0.00374907f
c145 12 Vss 0.0826302f
c146 10 Vss 0.0827668f
c147 6 Vss 0.00176834f
c148 4 Vss 0.0823731f
c149 2 Vss 0.0811326f
r150 95 104 1.16709
r151 95 96 0.470345
r152 93 102 0.326018
r153 92 100 0.551426
r154 92 93 4.16786
r155 91 100 0.551426
r156 90 91 13.3371
r157 86 100 0.0828784
r158 86 88 1.82344
r159 85 99 0.494161
r160 84 90 0.652036
r161 84 85 4.37625
r162 82 118 1.16709
r163 80 99 0.128424
r164 80 82 2.16729
r165 78 102 0.326018
r166 78 79 10.1279
r167 76 113 1.16709
r168 74 79 0.652036
r169 74 76 2.16729
r170 73 98 0.494161
r171 72 99 0.494161
r172 72 73 7.46046
r173 68 98 0.128424
r174 68 70 4.83471
r175 67 96 3.82922
r176 64 98 0.494161
r177 64 65 13.0037
r178 63 67 0.655813
r179 62 65 0.652036
r180 62 63 7.002
r181 49 118 0.197068
r182 46 49 1.2837
r183 42 113 0.197068
r184 42 44 1.2837
r185 38 46 0.0685365
r186 35 44 0.0685365
r187 31 104 0.0476429
r188 29 31 1.45875
r189 28 32 0.652036
r190 28 31 1.45875
r191 25 29 0.652036
r192 14 88 1.16709
r193 12 38 2.5674
r194 10 35 2.5674
r195 6 70 1.16709
r196 4 25 2.5674
r197 2 32 2.5674
.ends

.subckt PM_G3_DFFQ1_N1_CKN 2 6 8 18 28 33 50 Vss
c38 51 Vss 0.00127799f
c39 50 Vss 0.0053557f
c40 33 Vss 6.7412e-19
c41 28 Vss 0.00188103f
c42 18 Vss 8.89292e-19
c43 6 Vss 0.365937f
c44 2 Vss 0.00148239f
r45 50 51 14.6709
r46 46 51 0.652036
r47 33 50 0.531835
r48 28 46 4.00114
r49 18 33 1.16709
r50 8 18 6.4185
r51 6 18 6.4185
r52 2 28 1.16709
.ends

.subckt PM_G3_DFFQ1_N1_D 2 4 11 12 22 25 28 Vss
c27 28 Vss 0.00185315f
c28 25 Vss 4.49891e-19
c29 12 Vss 0.210787f
c30 11 Vss 2.35358e-19
c31 7 Vss 0.0247918f
c32 4 Vss 0.0830137f
c33 2 Vss 0.0713067f
r34 25 28 1.16709
r35 22 25 0.0364688
r36 15 28 0.0476429
r37 13 15 0.326018
r38 13 15 0.1167
r39 12 16 0.652036
r40 12 15 6.7686
r41 11 28 0.357321
r42 7 15 0.326018
r43 7 11 0.40845
r44 4 16 2.5674
r45 2 11 2.15895
.ends

.subckt PM_G3_DFFQ1_N1_X 2 4 8 17 20 23 35 39 41 47 Vss
c50 47 Vss 0.00138877f
c51 41 Vss 6.77172e-19
c52 39 Vss 0.0010541f
c53 35 Vss 0.00217231f
c54 23 Vss 7.53039e-20
c55 20 Vss 0.21062f
c56 17 Vss 0.0712602f
c57 15 Vss 0.0247918f
c58 8 Vss 0.0829593f
c59 2 Vss 0.00172036f
r60 44 47 1.16709
r61 41 44 2.08393
r62 37 39 4.33457
r63 36 41 0.0685365
r64 35 37 0.652036
r65 35 36 1.70882
r66 23 47 0.0476429
r67 21 23 0.326018
r68 21 23 0.1167
r69 20 24 0.652036
r70 20 23 6.7686
r71 17 47 0.357321
r72 15 23 0.326018
r73 15 17 0.40845
r74 8 24 2.5674
r75 4 17 2.15895
r76 2 39 1.16709
.ends

.subckt PM_G3_DFFQ1_N1_Q 2 16 Vss
c12 16 Vss 4.30842e-19
c13 2 Vss 0.00150258f
r14 16 19 0.0416786
r15 2 19 1.16709
.ends

.subckt G3_DFFQ1_N1  VSS CK VDD D Q
*
* Q	Q
* D	D
* VDD	VDD
* CK	CK
* VSS	VSS
XI1.X0 N_CKN_XI1.X0_D N_VDD_XI1.X0_PGD N_CK_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
XI2.X0 N_CKN_XI1.X0_D N_VSS_XI2.X0_PGD N_CK_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI5.X0 N_X_XI5.X0_D N_VSS_XI5.X0_PGD N_D_XI5.X0_CG N_CK_XI5.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI3.X0 N_Q_XI3.X0_D N_VDD_XI3.X0_PGD N_X_XI3.X0_CG N_CK_XI3.X0_PGS
+ N_VSS_XI3.X0_S TIGFET_HPNW1
XI4.X0 N_X_XI5.X0_D N_VDD_XI4.X0_PGD N_D_XI4.X0_CG N_CKN_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW1
XI0.X0 N_Q_XI3.X0_D N_VSS_XI0.X0_PGD N_X_XI0.X0_CG N_CKN_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW1
*
x_PM_G3_DFFQ1_N1_VSS N_VSS_XI1.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI5.X0_PGD N_VSS_XI3.X0_S N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_11_p
+ N_VSS_c_89_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_15_p N_VSS_c_3_p N_VSS_c_32_p
+ N_VSS_c_23_p N_VSS_c_33_p N_VSS_c_45_p N_VSS_c_20_p N_VSS_c_4_p N_VSS_c_34_p
+ N_VSS_c_16_p N_VSS_c_7_p N_VSS_c_22_p N_VSS_c_17_p N_VSS_c_85_p VSS
+ N_VSS_c_38_p N_VSS_c_29_p N_VSS_c_39_p N_VSS_c_48_p N_VSS_c_51_p N_VSS_c_52_p
+ N_VSS_c_30_p N_VSS_c_40_p N_VSS_c_53_p Vss PM_G3_DFFQ1_N1_VSS
x_PM_G3_DFFQ1_N1_CK N_CK_XI1.X0_CG N_CK_XI2.X0_CG N_CK_XI5.X0_PGS
+ N_CK_XI3.X0_PGS N_CK_c_122_n N_CK_c_123_n CK N_CK_c_129_p Vss
+ PM_G3_DFFQ1_N1_CK
x_PM_G3_DFFQ1_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI2.X0_S
+ N_VDD_XI3.X0_PGD N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_152_n N_VDD_c_250_p
+ N_VDD_c_153_n N_VDD_c_154_n N_VDD_c_155_n N_VDD_c_159_n N_VDD_c_163_n
+ N_VDD_c_164_n N_VDD_c_166_n N_VDD_c_172_n N_VDD_c_176_n N_VDD_c_182_n
+ N_VDD_c_183_n N_VDD_c_185_n N_VDD_c_188_n N_VDD_c_190_n N_VDD_c_195_n
+ N_VDD_c_199_n N_VDD_c_201_n N_VDD_c_203_n N_VDD_c_204_n N_VDD_c_205_n VDD
+ N_VDD_c_206_n N_VDD_c_208_n N_VDD_c_211_n Vss PM_G3_DFFQ1_N1_VDD
x_PM_G3_DFFQ1_N1_CKN N_CKN_XI1.X0_D N_CKN_XI4.X0_PGS N_CKN_XI0.X0_PGS
+ N_CKN_c_283_n N_CKN_c_268_n N_CKN_c_272_n N_CKN_c_274_n Vss PM_G3_DFFQ1_N1_CKN
x_PM_G3_DFFQ1_N1_D N_D_XI5.X0_CG N_D_XI4.X0_CG N_D_c_305_n N_D_c_306_n D
+ N_D_c_308_n N_D_c_312_n Vss PM_G3_DFFQ1_N1_D
x_PM_G3_DFFQ1_N1_X N_X_XI5.X0_D N_X_XI3.X0_CG N_X_XI0.X0_CG N_X_c_346_n
+ N_X_c_334_n N_X_c_354_n N_X_c_336_n N_X_c_337_n N_X_c_341_n N_X_c_343_n Vss
+ PM_G3_DFFQ1_N1_X
x_PM_G3_DFFQ1_N1_Q N_Q_XI3.X0_D Q Vss PM_G3_DFFQ1_N1_Q
cc_1 N_VSS_XI2.X0_PGS N_CK_XI5.X0_PGS 0.0029499f
cc_2 N_VSS_XI5.X0_PGD N_CK_XI5.X0_PGS 0.00158255f
cc_3 N_VSS_c_3_p N_CK_XI5.X0_PGS 8.20198e-19
cc_4 N_VSS_c_4_p N_CK_XI5.X0_PGS 4.62582e-19
cc_5 N_VSS_XI2.X0_PGD N_CK_c_122_n 4.16623e-19
cc_6 N_VSS_XI2.X0_PGS N_CK_c_123_n 4.26524e-19
cc_7 N_VSS_c_7_p CK 5.33707e-19
cc_8 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.00168612f
cc_9 N_VSS_XI0.X0_PGD N_VDD_XI3.X0_PGD 0.00189944f
cc_10 N_VSS_XI5.X0_PGD N_VDD_XI4.X0_PGD 0.00180681f
cc_11 N_VSS_c_11_p N_VDD_c_152_n 0.00168612f
cc_12 N_VSS_c_12_p N_VDD_c_153_n 0.00189944f
cc_13 N_VSS_c_13_p N_VDD_c_154_n 0.00180681f
cc_14 N_VSS_XI1.X0_S N_VDD_c_155_n 9.5668e-19
cc_15 N_VSS_c_15_p N_VDD_c_155_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_155_n 0.00321182f
cc_17 N_VSS_c_17_p N_VDD_c_155_n 0.00182807f
cc_18 N_VSS_c_15_p N_VDD_c_159_n 5.16845e-19
cc_19 N_VSS_c_3_p N_VDD_c_159_n 2.61925e-19
cc_20 N_VSS_c_20_p N_VDD_c_159_n 4.48125e-19
cc_21 N_VSS_c_7_p N_VDD_c_159_n 0.00922264f
cc_22 N_VSS_c_22_p N_VDD_c_163_n 0.00105444f
cc_23 N_VSS_c_23_p N_VDD_c_164_n 0.00239254f
cc_24 N_VSS_c_4_p N_VDD_c_164_n 9.55109e-19
cc_25 N_VSS_c_13_p N_VDD_c_166_n 2.43144e-19
cc_26 N_VSS_c_23_p N_VDD_c_166_n 0.00161703f
cc_27 N_VSS_c_4_p N_VDD_c_166_n 2.03837e-19
cc_28 N_VSS_c_7_p N_VDD_c_166_n 0.00131925f
cc_29 N_VSS_c_29_p N_VDD_c_166_n 0.00399563f
cc_30 N_VSS_c_30_p N_VDD_c_166_n 7.74609e-19
cc_31 N_VSS_c_3_p N_VDD_c_172_n 0.00179177f
cc_32 N_VSS_c_32_p N_VDD_c_172_n 3.92901e-19
cc_33 N_VSS_c_33_p N_VDD_c_172_n 8.51944e-19
cc_34 N_VSS_c_34_p N_VDD_c_172_n 3.99794e-19
cc_35 N_VSS_c_12_p N_VDD_c_176_n 3.37151e-19
cc_36 N_VSS_c_33_p N_VDD_c_176_n 0.00141228f
cc_37 N_VSS_c_34_p N_VDD_c_176_n 0.00112249f
cc_38 N_VSS_c_38_p N_VDD_c_176_n 0.00402042f
cc_39 N_VSS_c_39_p N_VDD_c_176_n 0.00326829f
cc_40 N_VSS_c_40_p N_VDD_c_176_n 7.74609e-19
cc_41 N_VSS_c_38_p N_VDD_c_182_n 0.00142104f
cc_42 N_VSS_c_23_p N_VDD_c_183_n 9.29543e-19
cc_43 N_VSS_c_4_p N_VDD_c_183_n 3.82294e-19
cc_44 N_VSS_XI4.X0_S N_VDD_c_185_n 3.7884e-19
cc_45 N_VSS_c_45_p N_VDD_c_185_n 4.73473e-19
cc_46 N_VSS_c_29_p N_VDD_c_185_n 0.00432522f
cc_47 N_VSS_c_45_p N_VDD_c_188_n 2.14355e-19
cc_48 N_VSS_c_48_p N_VDD_c_188_n 5.52785e-19
cc_49 N_VSS_XI4.X0_S N_VDD_c_190_n 9.5668e-19
cc_50 N_VSS_c_45_p N_VDD_c_190_n 0.00165395f
cc_51 N_VSS_c_51_p N_VDD_c_190_n 0.00302432f
cc_52 N_VSS_c_52_p N_VDD_c_190_n 0.00617602f
cc_53 N_VSS_c_53_p N_VDD_c_190_n 8.91588e-19
cc_54 N_VSS_c_33_p N_VDD_c_195_n 4.43871e-19
cc_55 N_VSS_c_34_p N_VDD_c_195_n 3.66936e-19
cc_56 N_VSS_c_39_p N_VDD_c_195_n 0.00106633f
cc_57 N_VSS_c_52_p N_VDD_c_195_n 0.00303537f
cc_58 N_VSS_c_3_p N_VDD_c_199_n 6.19689e-19
cc_59 N_VSS_c_20_p N_VDD_c_199_n 3.8721e-19
cc_60 N_VSS_c_15_p N_VDD_c_201_n 0.00303908f
cc_61 N_VSS_c_7_p N_VDD_c_201_n 2.94014e-19
cc_62 N_VSS_c_7_p N_VDD_c_203_n 0.00116322f
cc_63 N_VSS_c_29_p N_VDD_c_204_n 0.00102846f
cc_64 N_VSS_c_52_p N_VDD_c_205_n 0.00116512f
cc_65 N_VSS_c_3_p N_VDD_c_206_n 3.86162e-19
cc_66 N_VSS_c_20_p N_VDD_c_206_n 6.0892e-19
cc_67 N_VSS_c_3_p N_VDD_c_208_n 5.29489e-19
cc_68 N_VSS_c_33_p N_VDD_c_208_n 3.48267e-19
cc_69 N_VSS_c_34_p N_VDD_c_208_n 8.07896e-19
cc_70 N_VSS_c_23_p N_VDD_c_211_n 3.48267e-19
cc_71 N_VSS_c_4_p N_VDD_c_211_n 8.0279e-19
cc_72 N_VSS_XI1.X0_S N_CKN_XI1.X0_D 3.43419e-19
cc_73 N_VSS_c_15_p N_CKN_XI1.X0_D 3.48267e-19
cc_74 N_VSS_XI1.X0_S N_CKN_c_268_n 3.48267e-19
cc_75 N_VSS_c_15_p N_CKN_c_268_n 0.00105962f
cc_76 N_VSS_c_3_p N_CKN_c_268_n 7.53164e-19
cc_77 N_VSS_c_7_p N_CKN_c_268_n 5.38016e-19
cc_78 N_VSS_c_29_p N_CKN_c_272_n 2.21217e-19
cc_79 N_VSS_c_52_p N_CKN_c_272_n 0.00111539f
cc_80 N_VSS_c_3_p N_CKN_c_274_n 0.00220607f
cc_81 N_VSS_c_32_p N_CKN_c_274_n 8.60018e-19
cc_82 N_VSS_c_23_p N_CKN_c_274_n 2.36534e-19
cc_83 N_VSS_c_33_p N_CKN_c_274_n 7.62758e-19
cc_84 N_VSS_c_7_p N_CKN_c_274_n 0.00158805f
cc_85 N_VSS_c_85_p N_CKN_c_274_n 8.14378e-19
cc_86 N_VSS_c_38_p N_CKN_c_274_n 9.16986e-19
cc_87 N_VSS_c_29_p N_CKN_c_274_n 0.00110784f
cc_88 N_VSS_c_4_p N_D_XI5.X0_CG 0.00265616f
cc_89 N_VSS_c_89_p N_D_c_305_n 9.49637e-19
cc_90 N_VSS_XI5.X0_PGD N_D_c_306_n 3.8966e-19
cc_91 N_VSS_XI0.X0_PGD N_D_c_306_n 2.22031e-19
cc_92 N_VSS_c_3_p N_D_c_308_n 6.13924e-19
cc_93 N_VSS_c_23_p N_D_c_308_n 5.5494e-19
cc_94 N_VSS_c_20_p N_D_c_308_n 3.48267e-19
cc_95 N_VSS_c_4_p N_D_c_308_n 4.56568e-19
cc_96 N_VSS_c_3_p N_D_c_312_n 3.48267e-19
cc_97 N_VSS_c_23_p N_D_c_312_n 4.56568e-19
cc_98 N_VSS_c_20_p N_D_c_312_n 6.88619e-19
cc_99 N_VSS_c_4_p N_D_c_312_n 6.1245e-19
cc_100 N_VSS_XI4.X0_S N_X_XI5.X0_D 3.43419e-19
cc_101 N_VSS_c_45_p N_X_XI5.X0_D 3.48267e-19
cc_102 N_VSS_c_34_p N_X_XI0.X0_CG 0.00105235f
cc_103 N_VSS_XI5.X0_PGD N_X_c_334_n 2.09879e-19
cc_104 N_VSS_XI0.X0_PGD N_X_c_334_n 3.99472e-19
cc_105 N_VSS_c_38_p N_X_c_336_n 2.5064e-19
cc_106 N_VSS_XI4.X0_S N_X_c_337_n 3.48267e-19
cc_107 N_VSS_c_3_p N_X_c_337_n 4.71026e-19
cc_108 N_VSS_c_45_p N_X_c_337_n 5.69026e-19
cc_109 N_VSS_c_52_p N_X_c_337_n 2.04792e-19
cc_110 N_VSS_c_3_p N_X_c_341_n 0.00157847f
cc_111 N_VSS_c_52_p N_X_c_341_n 3.24972e-19
cc_112 N_VSS_c_3_p N_X_c_343_n 3.48267e-19
cc_113 N_VSS_c_4_p N_X_c_343_n 2.00604e-19
cc_114 N_VSS_XI3.X0_S N_Q_XI3.X0_D 3.43419e-19
cc_115 N_VSS_c_32_p N_Q_XI3.X0_D 3.48267e-19
cc_116 N_VSS_XI3.X0_S Q 3.48267e-19
cc_117 N_VSS_c_32_p Q 4.99861e-19
cc_118 N_CK_c_122_n N_VDD_XI1.X0_PGD 4.16623e-19
cc_119 N_CK_XI5.X0_PGS N_VDD_XI4.X0_PGD 2.40707e-19
cc_120 N_CK_c_123_n N_VDD_c_154_n 2.40707e-19
cc_121 CK N_VDD_c_155_n 5.04211e-19
cc_122 N_CK_c_129_p N_VDD_c_155_n 5.23418e-19
cc_123 N_CK_c_122_n N_VDD_c_159_n 0.00141086f
cc_124 CK N_VDD_c_159_n 0.00141439f
cc_125 N_CK_c_129_p N_VDD_c_159_n 0.00120361f
cc_126 N_CK_XI5.X0_PGS N_VDD_c_164_n 2.38687e-19
cc_127 N_CK_c_123_n N_VDD_c_164_n 5.38952e-19
cc_128 CK N_VDD_c_164_n 3.91916e-19
cc_129 N_CK_c_129_p N_VDD_c_164_n 2.80271e-19
cc_130 CK N_VDD_c_199_n 6.07878e-19
cc_131 N_CK_c_129_p N_VDD_c_199_n 4.67029e-19
cc_132 CK N_VDD_c_206_n 4.56568e-19
cc_133 N_CK_c_129_p N_VDD_c_206_n 0.00211811f
cc_134 N_CK_XI5.X0_PGS N_CKN_XI4.X0_PGS 4.11563e-19
cc_135 N_CK_XI5.X0_PGS N_CKN_c_283_n 2.73384e-19
cc_136 N_CK_XI5.X0_PGS N_D_XI5.X0_CG 4.28946e-19
cc_137 N_CK_XI5.X0_PGS N_D_XI4.X0_CG 2.59344e-19
cc_138 N_CK_XI5.X0_PGS N_D_c_312_n 0.00300565f
cc_139 N_CK_XI5.X0_PGS N_X_XI0.X0_CG 2.6404e-19
cc_140 N_CK_XI5.X0_PGS N_X_c_346_n 4.97357e-19
cc_141 N_CK_XI5.X0_PGS N_X_c_343_n 0.00630896f
cc_142 N_VDD_XI2.X0_S N_CKN_XI1.X0_D 3.43419e-19
cc_143 N_VDD_c_190_n N_CKN_XI4.X0_PGS 5.54393e-19
cc_144 N_VDD_c_190_n N_CKN_c_283_n 8.21431e-19
cc_145 N_VDD_XI2.X0_S N_CKN_c_268_n 3.48267e-19
cc_146 N_VDD_c_159_n N_CKN_c_268_n 5.01863e-19
cc_147 N_VDD_c_164_n N_CKN_c_268_n 5.35331e-19
cc_148 N_VDD_c_199_n N_CKN_c_268_n 6.42405e-19
cc_149 N_VDD_c_190_n N_CKN_c_272_n 7.71262e-19
cc_150 N_VDD_c_159_n N_CKN_c_274_n 4.68667e-19
cc_151 N_VDD_c_166_n N_CKN_c_274_n 3.15582e-19
cc_152 N_VDD_c_176_n N_CKN_c_274_n 4.71809e-19
cc_153 N_VDD_c_183_n N_CKN_c_274_n 2.56401e-19
cc_154 N_VDD_c_211_n N_D_XI4.X0_CG 0.00105644f
cc_155 N_VDD_XI3.X0_PGD N_D_c_306_n 2.08865e-19
cc_156 N_VDD_XI4.X0_PGD N_D_c_306_n 4.04053e-19
cc_157 N_VDD_XI2.X0_S N_X_XI5.X0_D 3.43419e-19
cc_158 N_VDD_c_164_n N_X_XI5.X0_D 3.48267e-19
cc_159 N_VDD_c_166_n N_X_XI5.X0_D 3.7884e-19
cc_160 N_VDD_c_208_n N_X_c_346_n 0.00269538f
cc_161 N_VDD_XI3.X0_PGD N_X_c_334_n 3.93054e-19
cc_162 N_VDD_XI4.X0_PGD N_X_c_334_n 2.22031e-19
cc_163 N_VDD_c_250_p N_X_c_354_n 8.95961e-19
cc_164 N_VDD_c_208_n N_X_c_354_n 2.97161e-19
cc_165 N_VDD_XI2.X0_S N_X_c_337_n 3.48267e-19
cc_166 N_VDD_c_164_n N_X_c_337_n 6.883e-19
cc_167 N_VDD_c_166_n N_X_c_337_n 5.3319e-19
cc_168 N_VDD_c_190_n N_X_c_337_n 8.74231e-19
cc_169 N_VDD_c_172_n N_X_c_341_n 6.5515e-19
cc_170 N_VDD_c_208_n N_X_c_341_n 4.80549e-19
cc_171 N_VDD_c_172_n N_X_c_343_n 4.85469e-19
cc_172 N_VDD_c_208_n N_X_c_343_n 6.1245e-19
cc_173 N_VDD_XI0.X0_S N_Q_XI3.X0_D 3.43419e-19
cc_174 N_VDD_c_176_n N_Q_XI3.X0_D 3.7884e-19
cc_175 N_VDD_c_188_n N_Q_XI3.X0_D 3.72199e-19
cc_176 N_VDD_XI0.X0_S Q 3.48267e-19
cc_177 N_VDD_c_176_n Q 5.12447e-19
cc_178 N_VDD_c_188_n Q 7.06537e-19
cc_179 N_CKN_XI4.X0_PGS N_D_XI4.X0_CG 0.00392964f
cc_180 N_CKN_XI4.X0_PGS N_X_c_334_n 0.00402435f
cc_181 N_CKN_c_283_n N_X_c_336_n 5.71169e-19
cc_182 N_CKN_c_274_n N_X_c_336_n 0.00120349f
cc_183 N_CKN_c_268_n N_X_c_337_n 2.66307e-19
cc_184 N_CKN_c_272_n N_X_c_337_n 8.08281e-19
cc_185 N_CKN_c_274_n N_X_c_337_n 6.2695e-19
cc_186 N_CKN_c_274_n N_X_c_341_n 7.98434e-19
cc_187 N_D_c_306_n N_X_c_334_n 0.00454934f
cc_188 N_D_c_306_n N_X_c_337_n 2.96904e-19
cc_189 N_D_c_308_n N_X_c_337_n 0.00151915f
cc_190 N_D_c_312_n N_X_c_337_n 9.22925e-19
cc_191 N_D_c_308_n N_X_c_341_n 0.00146206f
cc_192 N_D_c_312_n N_X_c_341_n 0.00103457f
cc_193 N_D_c_308_n N_X_c_343_n 4.56568e-19
cc_194 N_D_c_312_n N_X_c_343_n 0.00373298f
cc_195 N_X_c_336_n N_Q_XI3.X0_D 5.75967e-19
cc_196 N_X_c_336_n Q 8.57825e-19
*
.ends
*
*
.subckt DFFQ1_HPNW1 CK D Q VDD VSS
xgate (VSS CK VDD D Q) G3_DFFQ1_N1
.ends
*
* File: G1_INV1_N1.pex.netlist
* Created: Fri Feb 18 12:29:10 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G1_INV1_N1_VDD 2 5 15 28 30 34 37 43 Vss
c23 43 Vss 0.00628299f
c24 34 Vss 7.87399e-19
c25 30 Vss 0.00507852f
c26 28 Vss 0.00249774f
c27 26 Vss 0.00167323f
c28 15 Vss 0.0355813f
c29 14 Vss 0.102384f
c30 5 Vss 0.164813f
c31 2 Vss 0.00212755f
r32 34 43 1.16709
r33 32 34 2.45904
r34 31 37 0.326018
r35 30 32 0.652036
r36 30 31 7.41879
r37 26 37 0.326018
r38 26 28 5.08479
r39 17 43 0.214393
r40 15 17 1.4004
r41 14 18 0.652036
r42 14 17 1.5171
r43 11 15 0.652036
r44 5 18 2.5674
r45 5 11 2.5674
r46 2 28 1.16709
.ends

.subckt PM_G1_INV1_N1_A 2 4 9 12 22 25 28 Vss
c8 28 Vss 0.00718398f
c9 12 Vss 0.227852f
c10 9 Vss 0.0715834f
c11 7 Vss 0.0247918f
c12 4 Vss 0.0847975f
r13 25 28 1.16709
r14 22 25 0.0530455
r15 15 28 0.0476429
r16 13 15 0.326018
r17 13 15 0.1167
r18 12 16 0.652036
r19 12 15 6.7686
r20 9 28 0.357321
r21 7 15 0.326018
r22 7 9 0.40845
r23 4 16 2.5674
r24 2 9 2.15895
.ends

.subckt PM_G1_INV1_N1_VSS 3 6 14 27 32 37 49 50 56 Vss
c26 51 Vss 0.00126572f
c27 50 Vss 6.56738e-19
c28 49 Vss 0.00355297f
c29 37 Vss 0.0039192f
c30 32 Vss 0.00204286f
c31 27 Vss 6.63162e-19
c32 15 Vss 0.0358722f
c33 14 Vss 0.0994269f
c34 6 Vss 0.00276734f
c35 3 Vss 0.163777f
r36 51 56 0.326018
r37 49 56 0.326018
r38 49 50 7.46046
r39 45 50 0.652036
r40 32 51 5.08479
r41 27 37 1.16709
r42 27 45 2.41736
r43 17 37 0.238214
r44 15 17 1.45875
r45 14 18 0.652036
r46 14 17 1.45875
r47 11 15 0.652036
r48 6 32 1.16709
r49 3 18 2.5674
r50 3 11 2.5674
.ends

.subckt PM_G1_INV1_N1_Z 2 16 Vss
c11 2 Vss 0.00148239f
r12 16 19 0.125036
r13 2 19 1.16709
.ends

.subckt G1_INV1_N1  VDD A VSS Z
*
* Z	Z
* VSS	VSS
* A	A
* VDD	VDD
XI2.X0 N_Z_XI2.X0_D N_VSS_XI2.X0_PGD N_A_XI2.X0_CG N_VSS_XI2.X0_PGD
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI1.X0 N_Z_XI2.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW1
*
x_PM_G1_INV1_N1_VDD N_VDD_XI2.X0_S N_VDD_XI1.X0_PGD N_VDD_c_5_p N_VDD_c_4_p
+ N_VDD_c_6_p N_VDD_c_9_p VDD N_VDD_c_1_p Vss PM_G1_INV1_N1_VDD
x_PM_G1_INV1_N1_A N_A_XI2.X0_CG N_A_XI1.X0_CG N_A_c_29_p N_A_c_25_n A N_A_c_27_p
+ N_A_c_28_p Vss PM_G1_INV1_N1_A
x_PM_G1_INV1_N1_VSS N_VSS_XI2.X0_PGD N_VSS_XI1.X0_S N_VSS_c_34_n N_VSS_c_36_n
+ N_VSS_c_40_n N_VSS_c_42_n N_VSS_c_45_n N_VSS_c_46_n VSS Vss PM_G1_INV1_N1_VSS
x_PM_G1_INV1_N1_Z N_Z_XI2.X0_D Z Vss PM_G1_INV1_N1_Z
cc_1 N_VDD_c_1_p N_A_XI1.X0_CG 8.21222e-19
cc_2 N_VDD_XI1.X0_PGD N_A_c_25_n 4.26524e-19
cc_3 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00171093f
cc_4 N_VDD_c_4_p N_VSS_XI2.X0_PGD 4.197e-19
cc_5 N_VDD_c_5_p N_VSS_c_34_n 0.00171093f
cc_6 N_VDD_c_6_p N_VSS_c_34_n 4.82774e-19
cc_7 N_VDD_c_4_p N_VSS_c_36_n 0.00304634f
cc_8 N_VDD_c_6_p N_VSS_c_36_n 0.0015849f
cc_9 N_VDD_c_9_p N_VSS_c_36_n 9.51078e-19
cc_10 N_VDD_c_1_p N_VSS_c_36_n 3.5189e-19
cc_11 N_VDD_c_4_p N_VSS_c_40_n 3.08259e-19
cc_12 N_VDD_c_9_p N_VSS_c_40_n 0.00107037f
cc_13 N_VDD_c_4_p N_VSS_c_42_n 9.54992e-19
cc_14 N_VDD_c_9_p N_VSS_c_42_n 3.83199e-19
cc_15 N_VDD_c_1_p N_VSS_c_42_n 7.7548e-19
cc_16 N_VDD_c_6_p N_VSS_c_45_n 0.005791f
cc_17 N_VDD_c_6_p N_VSS_c_46_n 0.00172748f
cc_18 N_VDD_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_19 N_VDD_c_4_p N_Z_XI2.X0_D 3.48267e-19
cc_20 N_VDD_c_6_p N_Z_XI2.X0_D 3.55567e-19
cc_21 N_VDD_XI2.X0_S Z 3.48267e-19
cc_22 N_VDD_c_4_p Z 7.06424e-19
cc_23 N_VDD_c_6_p Z 4.789e-19
cc_24 N_A_c_25_n N_VSS_XI2.X0_PGD 4.21166e-19
cc_25 N_A_c_27_p N_VSS_c_36_n 0.00103813f
cc_26 N_A_c_28_p N_VSS_c_36_n 4.99367e-19
cc_27 N_A_c_29_p N_VSS_c_42_n 0.00250475f
cc_28 N_A_c_27_p N_VSS_c_42_n 4.99367e-19
cc_29 N_A_c_28_p N_VSS_c_42_n 0.0014909f
cc_30 N_VSS_XI1.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_31 N_VSS_c_40_n N_Z_XI2.X0_D 3.48267e-19
cc_32 N_VSS_XI1.X0_S Z 3.48267e-19
cc_33 N_VSS_c_40_n Z 7.85754e-19
cc_34 N_VSS_c_45_n Z 2.54816e-19
*
.ends
*
*
.subckt INV1_HPNW1 A Y VDD VSS
xgate (VDD A VSS Y) G1_INV1_N1
.ends
*
* File: G3_LATQ1_N1.pex.netlist
* Created: Tue Apr  5 11:43:13 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_LATQ1_N1_VDD 2 4 6 8 10 12 14 31 34 42 48 66 68 69 70 73 75 76 79
+ 81 85 89 91 92 94 100 105 Vss
c91 105 Vss 0.00462608f
c92 100 Vss 0.00538553f
c93 92 Vss 2.39889e-19
c94 91 Vss 3.56526e-19
c95 89 Vss 0.002537f
c96 87 Vss 0.00169593f
c97 85 Vss 9.25444e-19
c98 81 Vss 0.00432906f
c99 79 Vss 0.00113626f
c100 76 Vss 8.64506e-19
c101 75 Vss 0.00220359f
c102 73 Vss 0.00166444f
c103 70 Vss 8.63529e-19
c104 69 Vss 0.00558368f
c105 68 Vss 0.00685141f
c106 66 Vss 0.00204371f
c107 53 Vss 0.0307391f
c108 48 Vss 0.230209f
c109 42 Vss 0.0346914f
c110 41 Vss 0.0656875f
c111 34 Vss 6.95602e-20
c112 32 Vss 0.0348624f
c113 31 Vss 0.1003f
c114 14 Vss 0.0852073f
c115 12 Vss 0.00176834f
c116 10 Vss 0.0837105f
c117 8 Vss 0.0825478f
c118 6 Vss 0.0832227f
c119 4 Vss 0.0825437f
c120 2 Vss 0.00231819f
r121 87 94 0.326018
r122 87 89 4.83471
r123 85 105 1.16709
r124 83 85 2.16729
r125 82 92 0.494161
r126 81 94 0.326018
r127 81 82 7.41879
r128 79 100 1.16709
r129 77 92 0.128424
r130 77 79 2.16729
r131 75 92 0.494161
r132 75 76 4.41793
r133 71 91 0.0828784
r134 71 73 1.82344
r135 69 83 0.652036
r136 69 70 10.1279
r137 68 76 0.652036
r138 67 91 0.551426
r139 67 68 13.3371
r140 66 91 0.551426
r141 65 70 0.652036
r142 65 66 4.16786
r143 49 53 0.494161
r144 48 50 0.652036
r145 48 49 6.8853
r146 45 53 0.128424
r147 44 105 0.238214
r148 42 44 1.45875
r149 41 53 0.494161
r150 41 44 1.45875
r151 38 42 0.652036
r152 34 100 0.238214
r153 32 34 1.5171
r154 31 35 0.652036
r155 31 34 1.4004
r156 28 32 0.652036
r157 14 50 2.5674
r158 12 89 1.16709
r159 10 45 2.5674
r160 8 38 2.5674
r161 6 28 2.5674
r162 4 35 2.5674
r163 2 73 1.16709
.ends

.subckt PM_G3_LATQ1_N1_VSS 2 4 6 8 10 12 16 31 32 42 48 66 71 76 81 90 95 104
+ 106 107 108 113 114 119 129 130 132 Vss
c83 130 Vss 3.75522e-19
c84 129 Vss 4.28045e-19
c85 125 Vss 0.00127887f
c86 119 Vss 0.00326191f
c87 114 Vss 8.18866e-19
c88 113 Vss 0.00406272f
c89 108 Vss 8.24051e-19
c90 107 Vss 0.00164689f
c91 106 Vss 0.00145595f
c92 104 Vss 0.0042874f
c93 95 Vss 0.00390998f
c94 90 Vss 0.00430366f
c95 81 Vss 0.0025736f
c96 76 Vss 6.81193e-19
c97 71 Vss 9.80151e-19
c98 66 Vss 0.00132247f
c99 53 Vss 0.0307391f
c100 48 Vss 0.230436f
c101 42 Vss 0.0338877f
c102 41 Vss 0.0647949f
c103 32 Vss 0.0341879f
c104 31 Vss 0.0984533f
c105 16 Vss 0.085351f
c106 12 Vss 0.0838423f
c107 10 Vss 0.0825458f
c108 8 Vss 0.00178431f
c109 6 Vss 0.00237018f
c110 4 Vss 0.0842992f
c111 2 Vss 0.0825494f
r112 125 132 0.326018
r113 120 130 0.494161
r114 119 132 0.326018
r115 119 120 7.46046
r116 115 130 0.128424
r117 113 121 0.652036
r118 113 114 10.1279
r119 109 129 0.0828784
r120 107 130 0.494161
r121 107 108 4.37625
r122 106 114 0.652036
r123 105 129 0.551426
r124 105 106 4.16786
r125 104 129 0.551426
r126 103 108 0.652036
r127 103 104 13.3371
r128 81 125 4.83471
r129 76 95 1.16709
r130 76 121 2.16729
r131 71 90 1.16709
r132 71 115 2.16729
r133 66 109 1.82344
r134 49 53 0.494161
r135 48 50 0.652036
r136 48 49 6.8853
r137 45 53 0.128424
r138 44 95 0.238214
r139 42 44 1.45875
r140 41 53 0.494161
r141 41 44 1.45875
r142 38 42 0.652036
r143 34 90 0.238214
r144 32 34 1.45875
r145 31 35 0.652036
r146 31 34 1.45875
r147 28 32 0.652036
r148 16 50 2.5674
r149 12 45 2.5674
r150 10 38 2.5674
r151 8 81 1.16709
r152 6 66 1.16709
r153 4 28 2.5674
r154 2 35 2.5674
.ends

.subckt PM_G3_LATQ1_N1_G 2 4 6 14 15 22 31 37 Vss
c28 37 Vss 0.00243204f
c29 31 Vss 4.35685e-19
c30 29 Vss 0.0294543f
c31 22 Vss 0.152644f
c32 15 Vss 0.175771f
c33 14 Vss 3.53242e-19
c34 10 Vss 0.0247918f
c35 6 Vss 0.0835217f
c36 4 Vss 0.0840272f
c37 2 Vss 0.0715834f
r38 34 37 1.16709
r39 31 34 0.0833571
r40 23 29 0.494161
r41 22 24 0.652036
r42 22 23 4.84305
r43 19 29 0.128424
r44 18 37 0.0476429
r45 16 18 0.326018
r46 16 18 0.1167
r47 15 29 0.494161
r48 15 18 6.7686
r49 14 37 0.357321
r50 10 18 0.326018
r51 10 14 0.40845
r52 6 24 2.5674
r53 4 19 2.5674
r54 2 14 2.15895
.ends

.subckt PM_G3_LATQ1_N1_QN 2 4 6 8 17 20 23 40 45 48 53 69 Vss
c48 69 Vss 3.70906e-19
c49 53 Vss 0.0021144f
c50 48 Vss 0.00799496f
c51 45 Vss 0.00464908f
c52 40 Vss 7.75457e-19
c53 23 Vss 1.9003e-19
c54 20 Vss 0.213496f
c55 17 Vss 0.0714043f
c56 15 Vss 0.0247918f
c57 8 Vss 0.00402754f
c58 6 Vss 0.00402754f
c59 4 Vss 0.0829687f
r60 65 69 0.652036
r61 48 69 13.7956
r62 48 50 4.58464
r63 45 48 4.58464
r64 40 53 1.16709
r65 40 65 1.83386
r66 23 53 0.0476429
r67 21 23 0.326018
r68 21 23 0.1167
r69 20 24 0.652036
r70 20 23 6.7686
r71 17 53 0.357321
r72 15 23 0.326018
r73 15 17 0.40845
r74 8 50 1.16709
r75 6 45 1.16709
r76 4 24 2.5674
r77 2 17 2.15895
.ends

.subckt PM_G3_LATQ1_N1_GN 2 6 12 27 29 30 32 39 Vss
c46 39 Vss 0.00259221f
c47 32 Vss 2.5038e-19
c48 30 Vss 7.22041e-19
c49 29 Vss 0.00123575f
c50 27 Vss 9.12307e-19
c51 12 Vss 0.171268f
c52 6 Vss 0.17763f
c53 2 Vss 0.00172036f
r54 32 39 1.16709
r55 29 32 0.531835
r56 29 30 1.70882
r57 25 30 0.652036
r58 25 27 4.00114
r59 14 39 0.197068
r60 12 16 0.652036
r61 12 14 4.668
r62 6 16 5.835
r63 2 27 1.16709
.ends

.subckt PM_G3_LATQ1_N1_Q 2 18 Vss
c12 18 Vss 4.14768e-19
c13 2 Vss 0.00150258f
r14 2 18 1.16709
.ends

.subckt PM_G3_LATQ1_N1_D 2 4 10 14 Vss
c14 14 Vss 4.15825e-19
c15 10 Vss 1.35847e-19
c16 2 Vss 0.365962f
r17 14 17 0.0416786
r18 10 17 1.16709
r19 4 10 6.4185
r20 2 10 6.4185
.ends

.subckt G3_LATQ1_N1  VDD VSS G Q D
*
* D	D
* Q	Q
* G	G
* VSS	VSS
* VDD	VDD
XI2.X0 N_GN_XI2.X0_D N_VSS_XI2.X0_PGD N_G_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI0.X0 N_Q_XI0.X0_D N_VDD_XI0.X0_PGD N_QN_XI0.X0_CG N_VDD_XI0.X0_PGS
+ N_VSS_XI0.X0_S TIGFET_HPNW1
XI1.X0 N_GN_XI2.X0_D N_VDD_XI1.X0_PGD N_G_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
XI3.X0 N_Q_XI0.X0_D N_VSS_XI3.X0_PGD N_QN_XI3.X0_CG N_VSS_XI3.X0_PGS
+ N_VDD_XI3.X0_S TIGFET_HPNW1
XI5.X0 N_QN_XI5.X0_D N_VDD_XI5.X0_PGD N_D_XI5.X0_CG N_G_XI5.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
XI4.X0 N_QN_XI4.X0_D N_VSS_XI4.X0_PGD N_D_XI4.X0_CG N_GN_XI4.X0_PGS
+ N_VDD_XI3.X0_S TIGFET_HPNW1
*
x_PM_G3_LATQ1_N1_VDD N_VDD_XI2.X0_S N_VDD_XI0.X0_PGD N_VDD_XI0.X0_PGS
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI3.X0_S N_VDD_XI5.X0_PGD N_VDD_c_10_p
+ N_VDD_c_58_p N_VDD_c_7_p N_VDD_c_47_p N_VDD_c_16_p N_VDD_c_3_p N_VDD_c_8_p
+ N_VDD_c_38_p N_VDD_c_14_p N_VDD_c_15_p N_VDD_c_42_p N_VDD_c_20_p N_VDD_c_11_p
+ N_VDD_c_18_p N_VDD_c_5_p N_VDD_c_35_p N_VDD_c_41_p VDD N_VDD_c_23_p
+ N_VDD_c_19_p Vss PM_G3_LATQ1_N1_VDD
x_PM_G3_LATQ1_N1_VSS N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS N_VSS_XI0.X0_S
+ N_VSS_XI1.X0_S N_VSS_XI3.X0_PGD N_VSS_XI3.X0_PGS N_VSS_XI4.X0_PGD N_VSS_c_98_n
+ N_VSS_c_100_n N_VSS_c_101_n N_VSS_c_103_n N_VSS_c_104_n N_VSS_c_107_n
+ N_VSS_c_111_n N_VSS_c_115_n N_VSS_c_116_n N_VSS_c_120_n N_VSS_c_124_n
+ N_VSS_c_127_n N_VSS_c_128_n N_VSS_c_129_n N_VSS_c_130_n N_VSS_c_133_n
+ N_VSS_c_134_n N_VSS_c_135_n N_VSS_c_136_n VSS Vss PM_G3_LATQ1_N1_VSS
x_PM_G3_LATQ1_N1_G N_G_XI2.X0_CG N_G_XI1.X0_CG N_G_XI5.X0_PGS N_G_c_183_n
+ N_G_c_177_n N_G_c_179_n G N_G_c_181_n Vss PM_G3_LATQ1_N1_G
x_PM_G3_LATQ1_N1_QN N_QN_XI0.X0_CG N_QN_XI3.X0_CG N_QN_XI5.X0_D N_QN_XI4.X0_D
+ N_QN_c_205_n N_QN_c_206_n N_QN_c_208_n N_QN_c_210_n N_QN_c_213_n N_QN_c_215_n
+ N_QN_c_218_n N_QN_c_221_n Vss PM_G3_LATQ1_N1_QN
x_PM_G3_LATQ1_N1_GN N_GN_XI2.X0_D N_GN_XI4.X0_PGS N_GN_c_254_n N_GN_c_256_n
+ N_GN_c_279_n N_GN_c_285_n N_GN_c_260_n N_GN_c_262_n Vss PM_G3_LATQ1_N1_GN
x_PM_G3_LATQ1_N1_Q N_Q_XI0.X0_D Q Vss PM_G3_LATQ1_N1_Q
x_PM_G3_LATQ1_N1_D N_D_XI5.X0_CG N_D_XI4.X0_CG N_D_c_314_n D Vss
+ PM_G3_LATQ1_N1_D
cc_1 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00175469f
cc_2 N_VDD_XI0.X0_PGS N_VSS_XI2.X0_PGS 2.27468e-19
cc_3 N_VDD_c_3_p N_VSS_XI0.X0_S 9.5668e-19
cc_4 N_VDD_XI0.X0_PGD N_VSS_XI3.X0_PGD 0.00173629f
cc_5 N_VDD_c_5_p N_VSS_XI3.X0_PGS 2.46127e-19
cc_6 N_VDD_XI5.X0_PGD N_VSS_XI4.X0_PGD 2.27468e-19
cc_7 N_VDD_c_7_p N_VSS_c_98_n 0.00175469f
cc_8 N_VDD_c_8_p N_VSS_c_98_n 3.60588e-19
cc_9 N_VDD_c_8_p N_VSS_c_100_n 3.60588e-19
cc_10 N_VDD_c_10_p N_VSS_c_101_n 0.00173629f
cc_11 N_VDD_c_11_p N_VSS_c_101_n 2.60334e-19
cc_12 N_VDD_c_5_p N_VSS_c_103_n 7.75484e-19
cc_13 N_VDD_c_3_p N_VSS_c_104_n 0.00165395f
cc_14 N_VDD_c_14_p N_VSS_c_104_n 7.6714e-19
cc_15 N_VDD_c_15_p N_VSS_c_104_n 5.16845e-19
cc_16 N_VDD_c_16_p N_VSS_c_107_n 4.43871e-19
cc_17 N_VDD_c_8_p N_VSS_c_107_n 0.00161703f
cc_18 N_VDD_c_18_p N_VSS_c_107_n 9.31718e-19
cc_19 N_VDD_c_19_p N_VSS_c_107_n 3.48267e-19
cc_20 N_VDD_c_20_p N_VSS_c_111_n 9.36729e-19
cc_21 N_VDD_c_11_p N_VSS_c_111_n 0.00141228f
cc_22 N_VDD_c_5_p N_VSS_c_111_n 0.00291977f
cc_23 N_VDD_c_23_p N_VSS_c_111_n 3.5189e-19
cc_24 N_VDD_c_18_p N_VSS_c_115_n 0.00102583f
cc_25 N_VDD_c_16_p N_VSS_c_116_n 3.66936e-19
cc_26 N_VDD_c_8_p N_VSS_c_116_n 2.03837e-19
cc_27 N_VDD_c_18_p N_VSS_c_116_n 3.99794e-19
cc_28 N_VDD_c_19_p N_VSS_c_116_n 8.07896e-19
cc_29 N_VDD_c_20_p N_VSS_c_120_n 3.86045e-19
cc_30 N_VDD_c_11_p N_VSS_c_120_n 0.00112249f
cc_31 N_VDD_c_5_p N_VSS_c_120_n 9.54992e-19
cc_32 N_VDD_c_23_p N_VSS_c_120_n 8.1718e-19
cc_33 N_VDD_c_16_p N_VSS_c_124_n 0.00303537f
cc_34 N_VDD_c_3_p N_VSS_c_124_n 0.00544275f
cc_35 N_VDD_c_35_p N_VSS_c_124_n 0.00116512f
cc_36 N_VDD_c_3_p N_VSS_c_127_n 0.00305967f
cc_37 N_VDD_c_8_p N_VSS_c_128_n 0.00343927f
cc_38 N_VDD_c_38_p N_VSS_c_129_n 0.00106317f
cc_39 N_VDD_c_15_p N_VSS_c_130_n 0.00355199f
cc_40 N_VDD_c_11_p N_VSS_c_130_n 0.00567045f
cc_41 N_VDD_c_41_p N_VSS_c_130_n 9.48532e-19
cc_42 N_VDD_c_42_p N_VSS_c_133_n 0.00105938f
cc_43 N_VDD_c_8_p N_VSS_c_134_n 0.00557463f
cc_44 N_VDD_c_3_p N_VSS_c_135_n 8.91588e-19
cc_45 N_VDD_c_8_p N_VSS_c_136_n 7.74609e-19
cc_46 N_VDD_c_19_p N_G_XI1.X0_CG 8.09841e-19
cc_47 N_VDD_c_47_p N_G_XI5.X0_PGS 0.00162079f
cc_48 N_VDD_XI0.X0_PGD N_G_c_177_n 2.22031e-19
cc_49 N_VDD_XI1.X0_PGD N_G_c_177_n 3.93641e-19
cc_50 N_VDD_XI1.X0_PGS N_G_c_179_n 4.05198e-19
cc_51 N_VDD_c_3_p G 3.46645e-19
cc_52 N_VDD_c_3_p N_G_c_181_n 4.43544e-19
cc_53 N_VDD_XI3.X0_S N_QN_XI4.X0_D 3.43419e-19
cc_54 N_VDD_c_5_p N_QN_XI4.X0_D 3.48267e-19
cc_55 N_VDD_c_23_p N_QN_c_205_n 0.00269246f
cc_56 N_VDD_XI0.X0_PGD N_QN_c_206_n 4.05198e-19
cc_57 N_VDD_XI1.X0_PGD N_QN_c_206_n 2.0936e-19
cc_58 N_VDD_c_58_p N_QN_c_208_n 9.69462e-19
cc_59 N_VDD_c_23_p N_QN_c_208_n 2.60536e-19
cc_60 N_VDD_c_3_p N_QN_c_210_n 4.49462e-19
cc_61 N_VDD_c_20_p N_QN_c_210_n 4.57093e-19
cc_62 N_VDD_c_23_p N_QN_c_210_n 4.4444e-19
cc_63 N_VDD_XI3.X0_S N_QN_c_213_n 3.48267e-19
cc_64 N_VDD_c_5_p N_QN_c_213_n 9.00822e-19
cc_65 N_VDD_c_8_p N_QN_c_215_n 4.48879e-19
cc_66 N_VDD_c_11_p N_QN_c_215_n 3.93728e-19
cc_67 N_VDD_c_5_p N_QN_c_215_n 3.58217e-19
cc_68 N_VDD_c_3_p N_QN_c_218_n 6.61926e-19
cc_69 N_VDD_c_20_p N_QN_c_218_n 4.85469e-19
cc_70 N_VDD_c_23_p N_QN_c_218_n 6.1245e-19
cc_71 N_VDD_c_3_p N_QN_c_221_n 4.64547e-19
cc_72 N_VDD_XI2.X0_S N_GN_XI2.X0_D 3.43419e-19
cc_73 N_VDD_c_8_p N_GN_XI2.X0_D 3.7884e-19
cc_74 N_VDD_c_14_p N_GN_XI2.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_PGS N_GN_c_254_n 3.40151e-19
cc_76 N_VDD_c_47_p N_GN_c_254_n 3.20239e-19
cc_77 N_VDD_XI2.X0_S N_GN_c_256_n 3.48267e-19
cc_78 N_VDD_c_3_p N_GN_c_256_n 6.12365e-19
cc_79 N_VDD_c_8_p N_GN_c_256_n 5.32769e-19
cc_80 N_VDD_c_14_p N_GN_c_256_n 7.89245e-19
cc_81 N_VDD_c_18_p N_GN_c_260_n 2.2082e-19
cc_82 N_VDD_c_19_p N_GN_c_260_n 2.46105e-19
cc_83 N_VDD_c_18_p N_GN_c_262_n 2.68489e-19
cc_84 N_VDD_c_19_p N_GN_c_262_n 5.71759e-19
cc_85 N_VDD_XI3.X0_S N_Q_XI0.X0_D 3.43419e-19
cc_86 N_VDD_c_11_p N_Q_XI0.X0_D 3.7884e-19
cc_87 N_VDD_c_5_p N_Q_XI0.X0_D 3.48267e-19
cc_88 N_VDD_XI3.X0_S Q 3.48267e-19
cc_89 N_VDD_c_11_p Q 5.12447e-19
cc_90 N_VDD_c_5_p Q 7.06424e-19
cc_91 N_VDD_c_47_p N_D_XI5.X0_CG 4.07085e-19
cc_92 N_VSS_c_116_n N_G_XI2.X0_CG 0.00265616f
cc_93 N_VSS_c_116_n N_G_c_183_n 9.49637e-19
cc_94 N_VSS_XI2.X0_PGD N_G_c_177_n 3.99472e-19
cc_95 N_VSS_XI3.X0_PGD N_G_c_177_n 2.0936e-19
cc_96 N_VSS_c_107_n G 5.5494e-19
cc_97 N_VSS_c_116_n G 4.56568e-19
cc_98 N_VSS_c_124_n G 3.38887e-19
cc_99 N_VSS_c_107_n N_G_c_181_n 4.56568e-19
cc_100 N_VSS_c_116_n N_G_c_181_n 6.1245e-19
cc_101 N_VSS_c_120_n N_QN_XI3.X0_CG 8.05748e-19
cc_102 N_VSS_XI1.X0_S N_QN_XI5.X0_D 3.43419e-19
cc_103 N_VSS_c_115_n N_QN_XI5.X0_D 3.48267e-19
cc_104 N_VSS_XI2.X0_PGD N_QN_c_206_n 2.22031e-19
cc_105 N_VSS_XI3.X0_PGD N_QN_c_206_n 3.89061e-19
cc_106 N_VSS_c_130_n N_QN_c_210_n 2.91026e-19
cc_107 N_VSS_c_115_n N_QN_c_213_n 8.97415e-19
cc_108 N_VSS_c_111_n N_QN_c_215_n 3.5258e-19
cc_109 N_VSS_c_115_n N_QN_c_215_n 7.99552e-19
cc_110 N_VSS_c_130_n N_QN_c_215_n 6.85871e-19
cc_111 N_VSS_c_134_n N_QN_c_215_n 9.55516e-19
cc_112 N_VSS_c_107_n N_QN_c_221_n 5.43247e-19
cc_113 N_VSS_c_124_n N_QN_c_221_n 0.00168288f
cc_114 N_VSS_XI1.X0_S N_GN_XI2.X0_D 3.43419e-19
cc_115 N_VSS_c_115_n N_GN_XI2.X0_D 3.48267e-19
cc_116 N_VSS_c_103_n N_GN_XI4.X0_PGS 0.00163489f
cc_117 N_VSS_XI3.X0_PGS N_GN_c_254_n 6.77138e-19
cc_118 N_VSS_c_103_n N_GN_c_254_n 2.57527e-19
cc_119 N_VSS_XI1.X0_S N_GN_c_256_n 3.48267e-19
cc_120 N_VSS_c_115_n N_GN_c_256_n 4.97497e-19
cc_121 N_VSS_c_124_n N_GN_c_256_n 4.46497e-19
cc_122 N_VSS_c_120_n N_GN_c_260_n 2.46105e-19
cc_123 N_VSS_c_111_n N_GN_c_262_n 2.52506e-19
cc_124 N_VSS_c_120_n N_GN_c_262_n 5.99566e-19
cc_125 N_VSS_XI0.X0_S N_Q_XI0.X0_D 3.43419e-19
cc_126 N_VSS_c_104_n N_Q_XI0.X0_D 3.48267e-19
cc_127 N_VSS_XI0.X0_S Q 3.48267e-19
cc_128 N_VSS_c_104_n Q 7.78122e-19
cc_129 N_VSS_c_103_n N_D_XI5.X0_CG 4.07085e-19
cc_130 N_G_c_177_n N_QN_c_206_n 0.003965f
cc_131 G N_QN_c_210_n 5.07332e-19
cc_132 N_G_c_181_n N_QN_c_210_n 4.54925e-19
cc_133 N_G_c_181_n N_QN_c_218_n 0.00269321f
cc_134 N_G_c_179_n N_GN_c_254_n 0.00851239f
cc_135 N_G_c_177_n N_GN_c_256_n 3.2445e-19
cc_136 G N_GN_c_256_n 0.00153131f
cc_137 N_G_c_181_n N_GN_c_256_n 9.18093e-19
cc_138 N_G_c_177_n N_GN_c_279_n 3.7133e-19
cc_139 N_G_c_177_n N_GN_c_262_n 9.94034e-19
cc_140 N_G_c_181_n N_GN_c_262_n 2.41671e-19
cc_141 N_G_XI5.X0_PGS N_D_XI5.X0_CG 0.00409312f
cc_142 N_QN_c_206_n N_GN_XI4.X0_PGS 0.00182388f
cc_143 N_QN_c_213_n N_GN_c_256_n 7.80248e-19
cc_144 N_QN_c_215_n N_GN_c_279_n 8.96813e-19
cc_145 N_QN_c_215_n N_GN_c_285_n 0.00118168f
cc_146 N_QN_c_215_n N_GN_c_260_n 9.24681e-19
cc_147 N_QN_c_206_n N_GN_c_262_n 8.57779e-19
cc_148 N_QN_c_218_n N_GN_c_262_n 2.75519e-19
cc_149 N_QN_c_206_n N_D_XI5.X0_CG 3.26559e-19
cc_150 N_QN_c_213_n N_D_XI5.X0_CG 0.00101289f
cc_151 N_QN_c_213_n N_D_c_314_n 0.00127983f
cc_152 N_QN_c_213_n D 0.00141415f
cc_153 N_QN_c_215_n D 0.00146947f
cc_154 N_GN_c_285_n N_Q_XI0.X0_D 5.19956e-19
cc_155 N_GN_c_285_n Q 6.79271e-19
cc_156 N_GN_XI4.X0_PGS N_D_XI5.X0_CG 0.00503657f
cc_157 N_GN_c_254_n N_D_c_314_n 0.00333193f
cc_158 N_GN_c_260_n N_D_c_314_n 3.73302e-19
cc_159 N_GN_c_262_n N_D_c_314_n 8.5422e-19
cc_160 N_GN_c_260_n D 2.88184e-19
cc_161 N_GN_c_262_n D 3.48267e-19
*
.ends
*
*
.subckt LATQ1_HPNW1 D G Q VDD VSS
xgate (VDD VSS G Q D) G3_LATQ1_N1
.ends
*
* File: G4_MAJ3_N1.pex.netlist
* Created: Wed Mar  2 17:07:12 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MAJ3_N1_VDD 2 4 7 11 27 28 31 32 51 52 54 56 57 61 65 67 68 71 75
+ 78 79 80 90 95 Vss
c80 95 Vss 0.00471931f
c81 90 Vss 0.00455939f
c82 80 Vss 3.56526e-19
c83 79 Vss 3.56526e-19
c84 75 Vss 3.84406e-19
c85 71 Vss 9.33011e-19
c86 68 Vss 8.63529e-19
c87 67 Vss 0.00539264f
c88 65 Vss 0.00133146f
c89 61 Vss 0.00133512f
c90 57 Vss 0.00563423f
c91 56 Vss 0.0019972f
c92 54 Vss 0.00437281f
c93 52 Vss 0.00204371f
c94 51 Vss 8.63529e-19
c95 32 Vss 0.0336444f
c96 31 Vss 0.0988545f
c97 28 Vss 0.0346129f
c98 27 Vss 0.0990038f
c99 11 Vss 0.165071f
c100 7 Vss 0.165416f
c101 4 Vss 0.00207958f
c102 2 Vss 0.0026194f
r103 75 95 1.16709
r104 73 75 2.16729
r105 71 90 1.16709
r106 69 71 2.16729
r107 67 73 0.652036
r108 67 68 10.1279
r109 63 80 0.0828784
r110 63 65 1.82344
r111 59 79 0.0828784
r112 59 61 1.82344
r113 58 78 0.326018
r114 57 69 0.652036
r115 57 58 10.1279
r116 56 68 0.652036
r117 55 80 0.551426
r118 55 56 4.16786
r119 54 80 0.551426
r120 53 79 0.551426
r121 53 54 7.83557
r122 52 79 0.551426
r123 51 78 0.326018
r124 51 52 4.16786
r125 34 95 0.238214
r126 32 34 1.45875
r127 31 38 0.652036
r128 31 34 1.45875
r129 30 90 0.238214
r130 28 30 1.45875
r131 27 35 0.652036
r132 27 30 1.45875
r133 24 32 0.652036
r134 21 28 0.652036
r135 11 38 2.5674
r136 11 24 2.5674
r137 7 35 2.5674
r138 7 21 2.5674
r139 4 65 1.16709
r140 2 61 1.16709
.ends

.subckt PM_G4_MAJ3_N1_VSS 3 7 10 12 27 28 31 32 34 52 57 62 67 70 73 78 91 92 93
+ 94 95 104 114 115 117 Vss
c89 115 Vss 3.75522e-19
c90 114 Vss 3.75522e-19
c91 110 Vss 0.00127887f
c92 104 Vss 0.00344356f
c93 95 Vss 8.24051e-19
c94 94 Vss 0.00149351f
c95 93 Vss 8.24051e-19
c96 92 Vss 0.00149351f
c97 91 Vss 0.00617495f
c98 78 Vss 0.00390682f
c99 73 Vss 0.00498746f
c100 70 Vss 0.00347745f
c101 67 Vss 0.00294127f
c102 62 Vss 0.00184732f
c103 57 Vss 0.00132425f
c104 52 Vss 0.00115907f
c105 32 Vss 0.033157f
c106 31 Vss 0.0974849f
c107 28 Vss 0.0341879f
c108 27 Vss 0.0984533f
c109 12 Vss 0.00257143f
c110 10 Vss 0.00203161f
c111 7 Vss 0.166925f
c112 3 Vss 0.166819f
r113 110 117 0.326018
r114 106 115 0.494161
r115 105 114 0.494161
r116 104 117 0.326018
r117 104 105 7.46046
r118 100 115 0.128424
r119 96 114 0.128424
r120 94 115 0.494161
r121 94 95 4.37625
r122 92 114 0.494161
r123 92 93 4.37625
r124 91 95 0.652036
r125 90 93 0.652036
r126 90 91 18.8387
r127 70 106 8.04396
r128 67 70 5.41821
r129 62 110 4.83471
r130 57 78 1.16709
r131 57 100 2.16729
r132 52 73 1.16709
r133 52 96 2.16729
r134 34 78 0.238214
r135 32 34 1.45875
r136 31 38 0.652036
r137 31 34 1.45875
r138 30 73 0.238214
r139 28 30 1.45875
r140 27 35 0.652036
r141 27 30 1.45875
r142 24 32 0.652036
r143 21 28 0.652036
r144 12 67 1.16709
r145 10 62 1.16709
r146 7 38 2.5674
r147 7 24 2.5674
r148 3 35 2.5674
r149 3 21 2.5674
.ends

.subckt PM_G4_MAJ3_N1_A 2 4 6 8 11 15 29 32 53 57 69 72 74 77 79 81 82 85 87 90
+ 98 107 Vss
c80 110 Vss 1.14262e-19
c81 107 Vss 0.00533929f
c82 98 Vss 0.00481087f
c83 94 Vss 7.48717e-19
c84 87 Vss 6.11441e-19
c85 85 Vss 8.50217e-19
c86 82 Vss 4.65536e-19
c87 81 Vss 0.00274588f
c88 79 Vss 0.00488819f
c89 77 Vss 8.85587e-19
c90 74 Vss 0.00117147f
c91 73 Vss 0.00146569f
c92 72 Vss 0.00379017f
c93 69 Vss 0.00539132f
c94 57 Vss 0.135015f
c95 53 Vss 0.128028f
c96 32 Vss 0.2139f
c97 29 Vss 0.0749894f
c98 27 Vss 0.0247918f
c99 11 Vss 1.01176f
c100 8 Vss 0.00236553f
c101 6 Vss 0.00271742f
c102 4 Vss 0.0850321f
r103 107 110 0.1
r104 96 107 1.16709
r105 92 98 1.16709
r106 90 92 0.166714
r107 87 90 0.166714
r108 83 85 2.16729
r109 82 96 0.531835
r110 81 83 0.652036
r111 81 82 1.70882
r112 80 94 0.494161
r113 79 96 0.531835
r114 79 80 7.46046
r115 75 94 0.128424
r116 75 77 2.16729
r117 73 94 0.494161
r118 73 74 1.83386
r119 71 74 0.652036
r120 71 72 8.00229
r121 70 87 0.0685365
r122 69 72 0.652036
r123 69 70 10.2113
r124 55 57 4.53833
r125 52 110 0.262036
r126 52 53 2.26917
r127 49 52 2.26917
r128 44 57 0.00605528
r129 43 53 0.00605528
r130 40 55 0.00605528
r131 39 49 0.00605528
r132 35 98 0.0952857
r133 33 35 0.326018
r134 33 35 0.1167
r135 32 36 0.652036
r136 32 35 6.7686
r137 29 35 0.3335
r138 27 35 0.326018
r139 27 29 0.2334
r140 15 44 2.5674
r141 15 40 2.5674
r142 11 15 12.837
r143 11 43 2.5674
r144 11 15 12.837
r145 11 39 2.5674
r146 8 85 1.16709
r147 6 77 1.16709
r148 4 36 2.5674
r149 2 29 2.334
.ends

.subckt PM_G4_MAJ3_N1_BI 2 6 8 21 32 37 42 52 57 66 72 73 Vss
c61 73 Vss 3.33918e-19
c62 72 Vss 7.31231e-19
c63 66 Vss 0.00174781f
c64 57 Vss 0.00147766f
c65 52 Vss 0.00140496f
c66 42 Vss 0.0015273f
c67 37 Vss 0.00542097f
c68 32 Vss 0.00210957f
c69 21 Vss 0.0573997f
c70 6 Vss 0.0573997f
c71 2 Vss 0.0015046f
r72 72 73 0.65228
r73 71 72 3.42052
r74 66 71 0.65409
r75 42 57 1.16709
r76 42 73 2.1395
r77 37 52 1.16709
r78 37 77 12.0712
r79 37 66 1.96931
r80 32 49 1.16709
r81 32 77 2.08393
r82 21 57 0.50025
r83 18 52 0.50025
r84 8 21 1.80885
r85 6 18 1.80885
r86 2 49 0.1
.ends

.subckt PM_G4_MAJ3_N1_AI 2 7 11 31 37 46 51 60 69 Vss
c47 69 Vss 2.51637e-19
c48 60 Vss 0.00575758f
c49 51 Vss 0.00577434f
c50 46 Vss 9.64269e-19
c51 37 Vss 0.127837f
c52 36 Vss 1.23462e-19
c53 31 Vss 0.133405f
c54 7 Vss 1.0035f
c55 2 Vss 0.0015046f
r56 65 69 0.652036
r57 60 63 0.1
r58 51 63 1.16709
r59 51 69 13.7539
r60 46 65 2.16729
r61 36 60 0.262036
r62 36 37 2.334
r63 33 36 2.20433
r64 29 31 4.53833
r65 26 37 0.00605528
r66 25 31 0.00605528
r67 22 33 0.00605528
r68 21 29 0.00605528
r69 11 26 2.5674
r70 11 22 2.5674
r71 7 11 12.837
r72 7 25 2.5674
r73 7 11 12.837
r74 7 21 2.5674
r75 2 46 1.16709
.ends

.subckt PM_G4_MAJ3_N1_B 2 4 6 8 16 17 26 38 42 45 50 55 60 65 73 74 80 87 92 93
+ Vss
c73 93 Vss 4.59352e-19
c74 92 Vss 0.00214833f
c75 87 Vss 7.9499e-19
c76 80 Vss 8.69209e-19
c77 74 Vss 2.46868e-19
c78 73 Vss 0.00310209f
c79 65 Vss 0.00148695f
c80 60 Vss 0.00103393f
c81 55 Vss 0.004462f
c82 50 Vss 0.00190521f
c83 45 Vss 8.22554e-19
c84 38 Vss 0.00131454f
c85 26 Vss 0.0573997f
c86 20 Vss 0.0247918f
c87 17 Vss 0.0343999f
c88 16 Vss 0.183114f
c89 8 Vss 0.0573997f
c90 4 Vss 0.0714013f
c91 2 Vss 0.0847975f
r92 91 93 0.65228
r93 91 92 3.46076
r94 87 92 0.65228
r95 83 87 2.1006
r96 80 83 2.04225
r97 73 80 0.0685365
r98 73 74 10.3363
r99 69 74 0.652036
r100 50 65 1.16709
r101 50 93 2.1395
r102 45 60 1.16709
r103 45 83 0.0416786
r104 38 55 1.16709
r105 38 69 2.16729
r106 38 42 0.0833571
r107 36 55 0.0476429
r108 33 65 0.50025
r109 26 60 0.50025
r110 24 55 0.357321
r111 20 36 0.326018
r112 20 24 0.40845
r113 17 36 6.7686
r114 16 36 0.326018
r115 16 36 0.1167
r116 13 17 0.652036
r117 8 33 1.80885
r118 6 26 1.80885
r119 4 24 2.15895
r120 2 13 2.5674
.ends

.subckt PM_G4_MAJ3_N1_C 2 4 20 25 50 54 57 Vss
c27 57 Vss 0.00412628f
c28 54 Vss 7.72795e-19
c29 25 Vss 0.00139119f
c30 20 Vss 6.60907e-19
c31 4 Vss 0.00277614f
c32 2 Vss 0.00222834f
r33 50 57 1.08364
r34 50 54 9.25264
r35 25 57 0.521797
r36 20 54 0.521797
r37 4 25 1.16709
r38 2 20 1.16709
.ends

.subckt PM_G4_MAJ3_N1_Z 2 4 30 33 Vss
c33 30 Vss 0.00258707f
c34 4 Vss 0.00153036f
c35 2 Vss 0.00148239f
r36 33 35 4.50129
r37 30 33 4.668
r38 4 35 1.16709
r39 2 30 1.16709
.ends

.subckt G4_MAJ3_N1  VDD VSS A B C Z
*
* Z	Z
* C	C
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI6.X0 N_BI_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW1
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW1
XI5.X0 N_VSS_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_BI_XI6.X0_D TIGFET_HPNW1
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW1
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_BI_XI2.X0_CG N_AI_XI2.X0_PGD N_A_XI2.X0_S
+ TIGFET_HPNW1
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_B_XI4.X0_CG N_AI_XI4.X0_PGD N_C_XI4.X0_S
+ TIGFET_HPNW1
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_B_XI3.X0_CG N_A_XI3.X0_PGD N_A_XI3.X0_S
+ TIGFET_HPNW1
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_BI_XI1.X0_CG N_A_XI1.X0_PGD N_C_XI1.X0_S
+ TIGFET_HPNW1
*
x_PM_G4_MAJ3_N1_VDD N_VDD_XI6.X0_S N_VDD_XI8.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI7.X0_PGD N_VDD_c_65_p N_VDD_c_3_p N_VDD_c_66_p N_VDD_c_6_p
+ N_VDD_c_37_p N_VDD_c_9_p N_VDD_c_31_p N_VDD_c_13_p N_VDD_c_4_p N_VDD_c_36_p
+ N_VDD_c_38_p N_VDD_c_7_p N_VDD_c_40_p N_VDD_c_11_p N_VDD_c_15_p VDD
+ N_VDD_c_33_p N_VDD_c_34_p N_VDD_c_12_p N_VDD_c_16_p Vss PM_G4_MAJ3_N1_VDD
x_PM_G4_MAJ3_N1_VSS N_VSS_XI6.X0_PGD N_VSS_XI8.X0_PGD N_VSS_XI5.X0_D
+ N_VSS_XI7.X0_S N_VSS_c_83_n N_VSS_c_85_n N_VSS_c_86_n N_VSS_c_88_n
+ N_VSS_c_135_p N_VSS_c_89_n N_VSS_c_93_n N_VSS_c_97_n N_VSS_c_98_n
+ N_VSS_c_101_n N_VSS_c_102_n N_VSS_c_106_n N_VSS_c_110_n N_VSS_c_115_n
+ N_VSS_c_117_n N_VSS_c_118_n N_VSS_c_120_n N_VSS_c_121_n N_VSS_c_122_n
+ N_VSS_c_123_n VSS Vss PM_G4_MAJ3_N1_VSS
x_PM_G4_MAJ3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI2.X0_S N_A_XI3.X0_S
+ N_A_XI3.X0_PGD N_A_XI1.X0_PGD N_A_c_182_n N_A_c_171_n N_A_c_211_p N_A_c_213_p
+ N_A_c_172_n N_A_c_189_n N_A_c_177_n N_A_c_233_p N_A_c_199_p N_A_c_237_p
+ N_A_c_225_p N_A_c_236_p N_A_c_179_n A N_A_c_180_n N_A_c_207_p Vss
+ PM_G4_MAJ3_N1_A
x_PM_G4_MAJ3_N1_BI N_BI_XI6.X0_D N_BI_XI2.X0_CG N_BI_XI1.X0_CG N_BI_c_265_n
+ N_BI_c_253_n N_BI_c_262_n N_BI_c_269_n N_BI_c_270_n N_BI_c_271_n N_BI_c_273_n
+ N_BI_c_293_p N_BI_c_296_p Vss PM_G4_MAJ3_N1_BI
x_PM_G4_MAJ3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_315_n
+ N_AI_c_316_n N_AI_c_317_n N_AI_c_320_n N_AI_c_330_n N_AI_c_321_n Vss
+ PM_G4_MAJ3_N1_AI
x_PM_G4_MAJ3_N1_B N_B_XI6.X0_CG N_B_XI5.X0_CG N_B_XI4.X0_CG N_B_XI3.X0_CG
+ N_B_c_359_n N_B_c_377_n N_B_c_414_n N_B_c_361_n B N_B_c_380_n N_B_c_381_n
+ N_B_c_364_n N_B_c_386_n N_B_c_387_n N_B_c_371_n N_B_c_372_n N_B_c_405_n
+ N_B_c_408_n N_B_c_411_n N_B_c_412_n Vss PM_G4_MAJ3_N1_B
x_PM_G4_MAJ3_N1_C N_C_XI4.X0_S N_C_XI1.X0_S N_C_c_433_n N_C_c_435_n C
+ N_C_c_437_n N_C_c_436_n Vss PM_G4_MAJ3_N1_C
x_PM_G4_MAJ3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_463_n Z Vss PM_G4_MAJ3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017247f
cc_2 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172036f
cc_3 N_VDD_c_3_p N_VSS_c_83_n 0.0017247f
cc_4 N_VDD_c_4_p N_VSS_c_83_n 2.74208e-19
cc_5 N_VDD_c_4_p N_VSS_c_85_n 3.60588e-19
cc_6 N_VDD_c_6_p N_VSS_c_86_n 0.00172036f
cc_7 N_VDD_c_7_p N_VSS_c_86_n 2.46461e-19
cc_8 N_VDD_c_7_p N_VSS_c_88_n 3.60588e-19
cc_9 N_VDD_c_9_p N_VSS_c_89_n 4.43871e-19
cc_10 N_VDD_c_4_p N_VSS_c_89_n 0.00161703f
cc_11 N_VDD_c_11_p N_VSS_c_89_n 9.28314e-19
cc_12 N_VDD_c_12_p N_VSS_c_89_n 3.48267e-19
cc_13 N_VDD_c_13_p N_VSS_c_93_n 4.43871e-19
cc_14 N_VDD_c_7_p N_VSS_c_93_n 0.00161703f
cc_15 N_VDD_c_15_p N_VSS_c_93_n 8.31866e-19
cc_16 N_VDD_c_16_p N_VSS_c_93_n 3.48267e-19
cc_17 N_VDD_c_11_p N_VSS_c_97_n 8.49247e-19
cc_18 N_VDD_XI7.X0_PGD N_VSS_c_98_n 3.41313e-19
cc_19 N_VDD_c_15_p N_VSS_c_98_n 0.00507115f
cc_20 N_VDD_c_16_p N_VSS_c_98_n 9.58524e-19
cc_21 N_VDD_c_7_p N_VSS_c_101_n 0.00403287f
cc_22 N_VDD_c_9_p N_VSS_c_102_n 3.66936e-19
cc_23 N_VDD_c_4_p N_VSS_c_102_n 2.03837e-19
cc_24 N_VDD_c_11_p N_VSS_c_102_n 3.99794e-19
cc_25 N_VDD_c_12_p N_VSS_c_102_n 8.07896e-19
cc_26 N_VDD_c_13_p N_VSS_c_106_n 3.66936e-19
cc_27 N_VDD_c_7_p N_VSS_c_106_n 2.03837e-19
cc_28 N_VDD_c_15_p N_VSS_c_106_n 3.99794e-19
cc_29 N_VDD_c_16_p N_VSS_c_106_n 8.03027e-19
cc_30 N_VDD_c_9_p N_VSS_c_110_n 0.00303537f
cc_31 N_VDD_c_31_p N_VSS_c_110_n 0.00599011f
cc_32 N_VDD_c_13_p N_VSS_c_110_n 0.00284565f
cc_33 N_VDD_c_33_p N_VSS_c_110_n 0.00104624f
cc_34 N_VDD_c_34_p N_VSS_c_110_n 0.0010706f
cc_35 N_VDD_c_4_p N_VSS_c_115_n 0.00345066f
cc_36 N_VDD_c_36_p N_VSS_c_115_n 2.07484e-19
cc_37 N_VDD_c_37_p N_VSS_c_117_n 0.00106317f
cc_38 N_VDD_c_38_p N_VSS_c_118_n 2.07484e-19
cc_39 N_VDD_c_7_p N_VSS_c_118_n 0.00345066f
cc_40 N_VDD_c_40_p N_VSS_c_120_n 0.00106317f
cc_41 N_VDD_c_4_p N_VSS_c_121_n 0.00557569f
cc_42 N_VDD_c_4_p N_VSS_c_122_n 7.74609e-19
cc_43 N_VDD_c_7_p N_VSS_c_123_n 7.74609e-19
cc_44 N_VDD_c_16_p N_A_XI7.X0_CG 9.92565e-19
cc_45 N_VDD_XI7.X0_PGD N_A_c_171_n 3.90792e-19
cc_46 N_VDD_XI7.X0_PGD N_A_c_172_n 5.17967e-19
cc_47 N_VDD_c_4_p N_A_c_172_n 3.35498e-19
cc_48 N_VDD_c_7_p N_A_c_172_n 4.32724e-19
cc_49 N_VDD_c_15_p N_A_c_172_n 4.1682e-19
cc_50 N_VDD_c_16_p N_A_c_172_n 5.53168e-19
cc_51 N_VDD_c_11_p N_A_c_177_n 5.52801e-19
cc_52 N_VDD_c_12_p N_A_c_177_n 4.1541e-19
cc_53 N_VDD_c_31_p N_A_c_179_n 5.53687e-19
cc_54 N_VDD_c_31_p N_A_c_180_n 4.71537e-19
cc_55 N_VDD_XI6.X0_S N_BI_XI6.X0_D 3.43419e-19
cc_56 N_VDD_c_4_p N_BI_XI6.X0_D 3.70842e-19
cc_57 N_VDD_c_36_p N_BI_XI6.X0_D 3.72199e-19
cc_58 N_VDD_XI6.X0_S N_BI_c_253_n 3.48267e-19
cc_59 N_VDD_c_4_p N_BI_c_253_n 4.45573e-19
cc_60 N_VDD_c_36_p N_BI_c_253_n 5.2846e-19
cc_61 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_62 N_VDD_c_38_p N_AI_XI8.X0_D 3.72199e-19
cc_63 N_VDD_XI5.X0_PGD N_AI_XI2.X0_PGD 2.73831e-19
cc_64 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.86706e-19
cc_65 N_VDD_c_65_p N_AI_c_315_n 2.73831e-19
cc_66 N_VDD_c_66_p N_AI_c_316_n 2.86706e-19
cc_67 N_VDD_XI8.X0_S N_AI_c_317_n 3.48267e-19
cc_68 N_VDD_c_38_p N_AI_c_317_n 5.226e-19
cc_69 N_VDD_c_7_p N_AI_c_317_n 5.01863e-19
cc_70 N_VDD_c_15_p N_AI_c_320_n 0.00114922f
cc_71 N_VDD_c_7_p N_AI_c_321_n 2.39469e-19
cc_72 N_VDD_c_12_p N_B_XI5.X0_CG 0.00237871f
cc_73 N_VDD_XI5.X0_PGD N_B_c_359_n 3.9688e-19
cc_74 N_VDD_XI7.X0_PGD N_B_c_359_n 2.07132e-19
cc_75 N_VDD_c_31_p N_B_c_361_n 3.8625e-19
cc_76 N_VDD_c_11_p N_B_c_361_n 6.84022e-19
cc_77 N_VDD_c_12_p N_B_c_361_n 8.63725e-19
cc_78 N_VDD_c_11_p N_B_c_364_n 4.85469e-19
cc_79 N_VDD_c_12_p N_B_c_364_n 0.0014909f
cc_80 N_VDD_c_16_p N_B_c_364_n 5.33198e-19
cc_81 N_VSS_XI5.X0_D N_A_XI2.X0_S 3.43419e-19
cc_82 N_VSS_c_106_n N_A_c_182_n 0.00236445f
cc_83 N_VSS_XI8.X0_PGD N_A_c_171_n 3.86211e-19
cc_84 N_VSS_XI7.X0_S N_A_c_172_n 9.18655e-19
cc_85 N_VSS_c_97_n N_A_c_172_n 4.08476e-19
cc_86 N_VSS_c_98_n N_A_c_172_n 0.00149476f
cc_87 N_VSS_c_101_n N_A_c_172_n 2.91598e-19
cc_88 N_VSS_c_121_n N_A_c_172_n 2.51207e-19
cc_89 N_VSS_XI5.X0_D N_A_c_189_n 9.18655e-19
cc_90 N_VSS_c_97_n N_A_c_189_n 0.00202821f
cc_91 N_VSS_c_97_n N_A_c_177_n 0.0012307f
cc_92 N_VSS_c_135_p N_A_c_179_n 3.48564e-19
cc_93 N_VSS_c_93_n N_A_c_179_n 5.0102e-19
cc_94 N_VSS_c_106_n N_A_c_179_n 4.64764e-19
cc_95 N_VSS_c_110_n N_A_c_179_n 4.46304e-19
cc_96 N_VSS_c_93_n N_A_c_180_n 4.26083e-19
cc_97 N_VSS_c_102_n N_A_c_180_n 5.39888e-19
cc_98 N_VSS_c_106_n N_A_c_180_n 0.001324f
cc_99 N_VSS_XI5.X0_D N_BI_XI6.X0_D 3.43419e-19
cc_100 N_VSS_c_97_n N_BI_XI6.X0_D 3.48267e-19
cc_101 N_VSS_XI5.X0_D N_BI_c_253_n 3.48267e-19
cc_102 N_VSS_c_97_n N_BI_c_253_n 0.0010124f
cc_103 N_VSS_c_110_n N_BI_c_253_n 6.76595e-19
cc_104 N_VSS_c_121_n N_BI_c_253_n 6.07981e-19
cc_105 N_VSS_c_97_n N_BI_c_262_n 5.26238e-19
cc_106 N_VSS_c_121_n N_BI_c_262_n 7.0632e-19
cc_107 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_108 N_VSS_c_98_n N_AI_XI8.X0_D 3.48267e-19
cc_109 N_VSS_c_98_n N_AI_XI2.X0_PGD 2.04949e-19
cc_110 N_VSS_XI7.X0_S N_AI_c_317_n 3.48267e-19
cc_111 N_VSS_c_93_n N_AI_c_317_n 0.00173262f
cc_112 N_VSS_c_98_n N_AI_c_317_n 0.00129107f
cc_113 N_VSS_c_110_n N_AI_c_317_n 9.31051e-19
cc_114 N_VSS_c_98_n N_AI_c_320_n 0.00170897f
cc_115 N_VSS_c_98_n N_AI_c_330_n 2.82216e-19
cc_116 N_VSS_c_101_n N_AI_c_321_n 0.00934196f
cc_117 N_VSS_c_102_n N_B_XI6.X0_CG 9.70552e-19
cc_118 N_VSS_XI6.X0_PGD N_B_c_359_n 3.923e-19
cc_119 N_VSS_XI8.X0_PGD N_B_c_359_n 2.07132e-19
cc_120 N_VSS_c_110_n N_B_c_361_n 7.87668e-19
cc_121 N_VSS_c_97_n N_B_c_371_n 5.49592e-19
cc_122 N_VSS_c_101_n N_B_c_372_n 2.27662e-19
cc_123 N_VSS_XI7.X0_S N_C_XI4.X0_S 3.43419e-19
cc_124 N_VSS_c_98_n N_C_XI4.X0_S 3.48267e-19
cc_125 N_VSS_XI7.X0_S N_C_c_433_n 3.48267e-19
cc_126 N_VSS_c_98_n N_C_c_433_n 5.64614e-19
cc_127 N_A_c_199_p N_BI_XI2.X0_CG 2.16788e-19
cc_128 N_A_XI3.X0_PGD N_BI_c_265_n 8.79767e-19
cc_129 N_A_c_172_n N_BI_c_253_n 0.00115944f
cc_130 N_A_c_189_n N_BI_c_262_n 0.00163472f
cc_131 N_A_c_199_p N_BI_c_262_n 0.00112713f
cc_132 N_A_c_199_p N_BI_c_269_n 5.2034e-19
cc_133 N_A_c_189_n N_BI_c_270_n 3.37713e-19
cc_134 N_A_XI3.X0_PGD N_BI_c_271_n 0.00245019f
cc_135 N_A_c_207_p N_BI_c_271_n 3.56342e-19
cc_136 N_A_c_199_p N_BI_c_273_n 0.00124805f
cc_137 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174421f
cc_138 N_A_c_189_n N_AI_XI2.X0_PGD 8.48901e-19
cc_139 N_A_c_211_p N_AI_c_315_n 0.00195894f
cc_140 N_A_c_199_p N_AI_c_315_n 0.00178666f
cc_141 N_A_c_213_p N_AI_c_316_n 0.00202303f
cc_142 N_A_c_172_n N_AI_c_317_n 0.00165136f
cc_143 N_A_c_172_n N_AI_c_320_n 0.00201403f
cc_144 N_A_XI3.X0_PGD N_B_XI3.X0_CG 8.79767e-19
cc_145 N_A_c_207_p N_B_XI3.X0_CG 0.00234701f
cc_146 N_A_c_171_n N_B_c_359_n 0.0036024f
cc_147 N_A_c_172_n N_B_c_359_n 5.44634e-19
cc_148 N_A_c_180_n N_B_c_377_n 4.18059e-19
cc_149 N_A_c_172_n N_B_c_361_n 7.76373e-19
cc_150 N_A_c_189_n N_B_c_361_n 0.00128334f
cc_151 N_A_c_172_n N_B_c_380_n 3.26436e-19
cc_152 N_A_c_199_p N_B_c_381_n 3.96409e-19
cc_153 N_A_c_225_p N_B_c_381_n 9.9319e-19
cc_154 N_A_c_207_p N_B_c_381_n 4.87397e-19
cc_155 N_A_c_171_n N_B_c_364_n 3.81736e-19
cc_156 N_A_c_189_n N_B_c_364_n 5.63683e-19
cc_157 N_A_c_172_n N_B_c_386_n 3.8563e-19
cc_158 N_A_XI3.X0_PGD N_B_c_387_n 0.00312702f
cc_159 N_A_c_207_p N_B_c_387_n 0.00145837f
cc_160 N_A_c_189_n N_B_c_371_n 0.002414f
cc_161 N_A_c_233_p N_B_c_371_n 3.98537e-19
cc_162 N_A_c_199_p N_B_c_371_n 6.08993e-19
cc_163 N_A_c_172_n N_B_c_372_n 0.00197865f
cc_164 N_A_c_236_p N_C_c_435_n 2.22411e-19
cc_165 N_A_c_237_p N_C_c_436_n 4.03103e-19
cc_166 N_A_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_167 N_A_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_168 N_A_c_233_p N_Z_XI2.X0_D 3.48267e-19
cc_169 N_A_c_199_p N_Z_XI2.X0_D 9.18655e-19
cc_170 N_A_c_236_p N_Z_XI2.X0_D 3.48267e-19
cc_171 N_A_XI2.X0_S N_Z_c_463_n 3.48267e-19
cc_172 N_A_XI3.X0_S N_Z_c_463_n 3.48267e-19
cc_173 N_A_XI3.X0_PGD N_Z_c_463_n 5.57521e-19
cc_174 N_A_c_189_n N_Z_c_463_n 9.24e-19
cc_175 N_A_c_233_p N_Z_c_463_n 7.8992e-19
cc_176 N_A_c_199_p N_Z_c_463_n 0.00158543f
cc_177 N_A_c_236_p N_Z_c_463_n 8.08848e-19
cc_178 N_BI_XI2.X0_CG N_AI_XI2.X0_PGD 8.63152e-19
cc_179 N_BI_c_270_n N_AI_XI2.X0_PGD 0.00312702f
cc_180 N_BI_c_253_n N_AI_c_317_n 3.22835e-19
cc_181 N_BI_c_262_n N_AI_c_320_n 3.68388e-19
cc_182 N_BI_c_270_n N_AI_c_330_n 2.00604e-19
cc_183 N_BI_c_262_n N_B_c_361_n 0.00136623f
cc_184 N_BI_c_262_n N_B_c_380_n 6.77523e-19
cc_185 N_BI_c_270_n N_B_c_380_n 4.99367e-19
cc_186 N_BI_c_269_n N_B_c_381_n 0.00186236f
cc_187 N_BI_c_271_n N_B_c_381_n 4.99367e-19
cc_188 N_BI_c_273_n N_B_c_381_n 0.00166575f
cc_189 N_BI_c_270_n N_B_c_386_n 0.00513784f
cc_190 N_BI_c_271_n N_B_c_386_n 7.2092e-19
cc_191 N_BI_c_269_n N_B_c_387_n 4.99367e-19
cc_192 N_BI_c_270_n N_B_c_387_n 6.22265e-19
cc_193 N_BI_c_271_n N_B_c_387_n 0.00499463f
cc_194 N_BI_c_262_n N_B_c_371_n 0.00525284f
cc_195 N_BI_c_262_n N_B_c_405_n 2.67017e-19
cc_196 N_BI_c_273_n N_B_c_405_n 0.0013533f
cc_197 N_BI_c_293_p N_B_c_405_n 0.00340518f
cc_198 N_BI_c_262_n N_B_c_408_n 4.99817e-19
cc_199 N_BI_c_273_n N_B_c_408_n 9.35879e-19
cc_200 N_BI_c_296_p N_B_c_408_n 7.59935e-19
cc_201 N_BI_c_293_p N_B_c_411_n 0.00181541f
cc_202 N_BI_c_262_n N_B_c_412_n 0.00138818f
cc_203 N_BI_c_273_n N_B_c_412_n 8.23093e-19
cc_204 N_BI_c_262_n N_C_c_437_n 3.43796e-19
cc_205 N_BI_c_262_n N_C_c_436_n 7.49861e-19
cc_206 N_BI_c_269_n N_C_c_436_n 9.95458e-19
cc_207 N_BI_c_296_p N_C_c_436_n 3.37189e-19
cc_208 N_BI_c_262_n N_Z_c_463_n 0.00187303f
cc_209 N_BI_c_269_n N_Z_c_463_n 0.00192908f
cc_210 N_BI_c_270_n N_Z_c_463_n 8.66889e-19
cc_211 N_BI_c_271_n N_Z_c_463_n 8.66889e-19
cc_212 N_BI_c_273_n N_Z_c_463_n 7.39431e-19
cc_213 N_BI_c_293_p N_Z_c_463_n 0.00210701f
cc_214 N_BI_c_296_p N_Z_c_463_n 9.92397e-19
cc_215 N_AI_XI2.X0_PGD N_B_c_414_n 8.79767e-19
cc_216 N_AI_c_330_n N_B_c_414_n 0.00234701f
cc_217 N_AI_c_320_n N_B_c_380_n 5.22873e-19
cc_218 N_AI_c_330_n N_B_c_380_n 4.87397e-19
cc_219 N_AI_XI2.X0_PGD N_B_c_386_n 0.00312702f
cc_220 N_AI_c_320_n N_B_c_386_n 4.3265e-19
cc_221 N_AI_c_330_n N_B_c_386_n 0.00145837f
cc_222 N_AI_c_320_n N_B_c_372_n 0.00441104f
cc_223 N_AI_c_320_n N_B_c_405_n 3.85994e-19
cc_224 N_AI_c_320_n N_C_c_433_n 0.00187508f
cc_225 N_AI_c_317_n N_C_c_437_n 2.87718e-19
cc_226 N_AI_c_320_n N_C_c_437_n 8.98954e-19
cc_227 N_AI_c_320_n N_C_c_436_n 5.19511e-19
cc_228 N_AI_XI2.X0_PGD N_Z_c_463_n 2.98914e-19
cc_229 N_B_c_371_n N_C_c_433_n 8.83421e-19
cc_230 N_B_c_381_n N_C_c_436_n 9.42245e-19
cc_231 N_B_c_371_n N_C_c_436_n 2.24447e-19
cc_232 N_B_c_408_n N_C_c_436_n 0.00527131f
cc_233 N_B_c_380_n N_Z_c_463_n 0.00210511f
cc_234 N_B_c_381_n N_Z_c_463_n 0.00187303f
cc_235 N_B_c_387_n N_Z_c_463_n 8.66889e-19
cc_236 N_B_c_405_n N_Z_c_463_n 4.75654e-19
cc_237 N_C_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_238 N_C_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_239 N_C_c_433_n N_Z_XI4.X0_D 3.48267e-19
cc_240 N_C_c_435_n N_Z_XI4.X0_D 3.48267e-19
cc_241 N_C_XI4.X0_S N_Z_c_463_n 3.48267e-19
cc_242 N_C_XI1.X0_S N_Z_c_463_n 3.48267e-19
cc_243 N_C_c_433_n N_Z_c_463_n 5.74266e-19
cc_244 N_C_c_435_n N_Z_c_463_n 5.79289e-19
cc_245 N_C_c_436_n N_Z_c_463_n 4.30842e-19
*
.ends
*
*
.subckt MAJ3_HPNW1 A B C Y VDD VSS
xgate (VDD VSS A B C Y) G4_MAJ3_N1
.ends
*
* File: G3_MIN3_T6_N1.pex.netlist
* Created: Sun Apr 10 19:28:11 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MIN3_T6_N1_VSS 2 4 6 10 12 22 27 32 37 40 42 45 60 65 70 75 88 89
+ 93 99 102 103 108 Vss
c79 109 Vss 6.38121e-19
c80 108 Vss 0.00185802f
c81 103 Vss 0.00201533f
c82 99 Vss 0.0091126f
c83 94 Vss 0.00136513f
c84 93 Vss 0.00679427f
c85 89 Vss 6.52641e-19
c86 88 Vss 0.00390198f
c87 75 Vss 0.00302736f
c88 70 Vss 3.56438e-22
c89 65 Vss 0.00159414f
c90 60 Vss 9.05888e-19
c91 45 Vss 0.0850774f
c92 42 Vss 0.0849587f
c93 37 Vss 0.0679309f
c94 32 Vss 0.103393f
c95 27 Vss 0.306892f
c96 22 Vss 0.138043f
c97 12 Vss 0.00262003f
c98 10 Vss 0.0805405f
c99 6 Vss 0.0807339f
c100 4 Vss 0.00185192f
c101 2 Vss 0.0794633f
r102 107 108 3.66771
r103 103 107 0.655813
r104 100 109 0.494161
r105 100 102 12.1285
r106 99 108 0.652036
r107 99 102 0.87525
r108 95 109 0.128424
r109 93 109 0.494161
r110 93 94 10.0862
r111 88 94 0.652036
r112 87 89 0.655813
r113 87 88 9.08593
r114 70 103 1.82344
r115 65 95 4.33457
r116 60 75 1.16709
r117 60 89 1.82344
r118 45 47 1.8672
r119 42 44 1.8672
r120 40 75 0.50025
r121 37 40 1.92555
r122 33 47 0.0685365
r123 32 34 0.652036
r124 32 33 2.8008
r125 29 47 0.5835
r126 28 42 0.0685365
r127 27 45 0.0685365
r128 27 28 10.9698
r129 24 44 0.5835
r130 23 37 0.0685365
r131 22 44 0.0685365
r132 22 23 4.7847
r133 12 70 1.16709
r134 10 34 2.5674
r135 6 29 2.5674
r136 4 65 1.16709
r137 2 24 2.5674
.ends

.subckt PM_G3_MIN3_T6_N1_VDD 2 4 8 10 12 22 27 32 42 45 60 61 63 65 69 71 73 78
+ 81 83 Vss
c82 83 Vss 0.00427875f
c83 79 Vss 7.70868e-19
c84 78 Vss 0.00350656f
c85 73 Vss 0.00126506f
c86 71 Vss 0.0122742f
c87 69 Vss 0.00176475f
c88 65 Vss 0.00137661f
c89 63 Vss 7.01183e-19
c90 62 Vss 0.00177567f
c91 61 Vss 0.00769188f
c92 60 Vss 0.00512434f
c93 45 Vss 0.0848894f
c94 42 Vss 0.0854608f
c95 38 Vss 0.0711342f
c96 32 Vss 0.106688f
c97 27 Vss 0.309245f
c98 22 Vss 0.14138f
c99 12 Vss 0.0779484f
c100 10 Vss 0.0024321f
c101 8 Vss 0.0787627f
c102 4 Vss 0.0785563f
c103 2 Vss 0.00185192f
r104 78 81 0.349767
r105 77 78 3.66771
r106 73 81 0.306046
r107 73 75 1.82344
r108 72 79 0.494161
r109 71 77 0.652036
r110 71 72 13.0037
r111 67 79 0.128424
r112 67 69 4.33457
r113 65 83 1.16709
r114 63 65 1.82344
r115 61 79 0.494161
r116 61 62 10.0862
r117 60 63 0.655813
r118 59 62 0.652036
r119 59 60 9.08593
r120 45 46 1.8672
r121 42 43 1.8672
r122 38 83 0.50025
r123 38 40 1.92555
r124 33 45 0.0685365
r125 32 34 0.652036
r126 32 33 2.8008
r127 29 45 0.5835
r128 28 43 0.0685365
r129 27 46 0.0685365
r130 27 28 10.9698
r131 24 42 0.5835
r132 23 40 0.0685365
r133 22 42 0.0685365
r134 22 23 4.7847
r135 12 34 2.5674
r136 10 75 1.16709
r137 8 29 2.5674
r138 4 24 2.5674
r139 2 69 1.16709
.ends

.subckt PM_G3_MIN3_T6_N1_Z 2 4 6 8 48 56 59 61 Vss
c50 61 Vss 0.00482259f
c51 56 Vss 0.00183713f
c52 48 Vss 0.00151912f
c53 8 Vss 0.00176753f
c54 6 Vss 0.00171956f
c55 4 Vss 6.64706e-19
c56 2 Vss 6.16734e-19
r57 61 63 2.79246
r58 59 61 0.125036
r59 56 59 2.50071
r60 51 61 10.7364
r61 51 53 2.79246
r62 48 51 2.62575
r63 8 63 1.16709
r64 6 56 1.16709
r65 4 53 1.16709
r66 2 48 1.16709
.ends

.subckt PM_G3_MIN3_T6_N1_C 2 4 6 8 14 20 29 32 37 42 Vss
c31 42 Vss 0.0053281f
c32 37 Vss 0.00169525f
c33 32 Vss 0.00511278f
c34 29 Vss 5.02822e-19
c35 20 Vss 0.268178f
c36 14 Vss 0.269305f
r37 32 42 1.16709
r38 29 37 1.16709
r39 29 32 10.0654
r40 20 42 0.50025
r41 14 37 0.50025
r42 6 8 7.5855
r43 6 20 1.80885
r44 2 4 7.5855
r45 2 14 1.80885
.ends

.subckt PM_G3_MIN3_T6_N1_B 2 4 6 8 17 18 26 32 35 Vss
c28 35 Vss 0.00171406f
c29 32 Vss 3.1388e-19
c30 26 Vss 0.0844898f
c31 18 Vss 0.0345851f
c32 17 Vss 0.0963137f
c33 6 Vss 0.292132f
c34 2 Vss 0.340186f
r35 29 35 1.16709
r36 29 32 0.0729375
r37 24 35 0.0476429
r38 24 26 1.92555
r39 17 19 0.652036
r40 17 18 2.8008
r41 14 26 0.0685365
r42 13 18 0.652036
r43 6 8 7.5855
r44 6 19 2.5674
r45 4 14 2.5674
r46 2 4 7.5855
r47 2 13 2.5674
.ends

.subckt PM_G3_MIN3_T6_N1_A 2 4 6 8 29 34 37 41 46 Vss
c28 46 Vss 0.00547458f
c29 41 Vss 0.00144837f
c30 37 Vss 0.00108816f
c31 34 Vss 5.02933e-19
c32 29 Vss 3.18404e-19
c33 26 Vss 0.087104f
c34 6 Vss 0.296947f
c35 2 Vss 0.267858f
r36 37 46 1.16709
r37 34 37 0.0833571
r38 29 41 1.16709
r39 29 37 5.03269
r40 24 46 0.0476429
r41 24 26 1.92555
r42 19 26 0.0685365
r43 17 41 0.50025
r44 8 19 2.5674
r45 6 8 7.5855
r46 4 17 1.80885
r47 2 4 7.5855
.ends

.subckt G3_MIN3_T6_N1  VSS VDD Z C B A
*
* A	A
* B	B
* C	C
* Z	Z
* VDD	VDD
* VSS	VSS
XI9.X0 N_Z_XI9.X0_D N_VSS_XI9.X0_PGD N_C_XI9.X0_CG N_B_XI9.X0_PGS N_VDD_XI9.X0_S
+ TIGFET_HPNW1
XI6.X0 N_Z_XI6.X0_D N_VDD_XI6.X0_PGD N_C_XI6.X0_CG N_B_XI6.X0_PGS N_VSS_XI6.X0_S
+ TIGFET_HPNW1
XI11.X0 N_Z_XI11.X0_D N_VSS_XI11.X0_PGD N_A_XI11.X0_CG N_B_XI11.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW1
XI10.X0 N_Z_XI10.X0_D N_VDD_XI10.X0_PGD N_A_XI10.X0_CG N_B_XI10.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW1
XI8.X0 N_Z_XI11.X0_D N_VSS_XI8.X0_PGD N_C_XI8.X0_CG N_A_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW1
XI7.X0 N_Z_XI10.X0_D N_VDD_XI7.X0_PGD N_C_XI7.X0_CG N_A_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW1
*
x_PM_G3_MIN3_T6_N1_VSS N_VSS_XI9.X0_PGD N_VSS_XI6.X0_S N_VSS_XI11.X0_PGD
+ N_VSS_XI8.X0_PGD N_VSS_XI7.X0_S N_VSS_c_8_p N_VSS_c_24_p N_VSS_c_27_p
+ N_VSS_c_9_p N_VSS_c_15_p N_VSS_c_16_p N_VSS_c_61_p N_VSS_c_10_p N_VSS_c_2_p
+ N_VSS_c_6_p N_VSS_c_11_p N_VSS_c_12_p N_VSS_c_13_p N_VSS_c_19_p N_VSS_c_28_p
+ VSS N_VSS_c_31_p N_VSS_c_76_p Vss PM_G3_MIN3_T6_N1_VSS
x_PM_G3_MIN3_T6_N1_VDD N_VDD_XI9.X0_S N_VDD_XI6.X0_PGD N_VDD_XI10.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI7.X0_PGD N_VDD_c_87_n N_VDD_c_150_p N_VDD_c_160_p
+ N_VDD_c_153_p N_VDD_c_152_p N_VDD_c_88_n N_VDD_c_93_n N_VDD_c_99_n
+ N_VDD_c_100_n N_VDD_c_102_n N_VDD_c_105_n N_VDD_c_108_n N_VDD_c_142_p VDD
+ N_VDD_c_111_n Vss PM_G3_MIN3_T6_N1_VDD
x_PM_G3_MIN3_T6_N1_Z N_Z_XI9.X0_D N_Z_XI6.X0_D N_Z_XI11.X0_D N_Z_XI10.X0_D
+ N_Z_c_170_n N_Z_c_176_n Z N_Z_c_180_n Vss PM_G3_MIN3_T6_N1_Z
x_PM_G3_MIN3_T6_N1_C N_C_XI9.X0_CG N_C_XI6.X0_CG N_C_XI8.X0_CG N_C_XI7.X0_CG
+ N_C_c_212_n N_C_c_213_n C N_C_c_214_n N_C_c_215_n N_C_c_216_n Vss
+ PM_G3_MIN3_T6_N1_C
x_PM_G3_MIN3_T6_N1_B N_B_XI9.X0_PGS N_B_XI6.X0_PGS N_B_XI11.X0_PGS
+ N_B_XI10.X0_PGS N_B_c_247_n N_B_c_248_n N_B_c_256_n B N_B_c_258_n Vss
+ PM_G3_MIN3_T6_N1_B
x_PM_G3_MIN3_T6_N1_A N_A_XI11.X0_CG N_A_XI10.X0_CG N_A_XI8.X0_PGS N_A_XI7.X0_PGS
+ N_A_c_272_n A N_A_c_276_n N_A_c_282_n N_A_c_283_n Vss PM_G3_MIN3_T6_N1_A
cc_1 N_VSS_XI6.X0_S N_VDD_XI9.X0_S 4.21365e-19
cc_2 N_VSS_c_2_p N_VDD_XI9.X0_S 3.8999e-19
cc_3 N_VSS_XI9.X0_PGD N_VDD_XI6.X0_PGD 6.1888e-19
cc_4 N_VSS_XI11.X0_PGD N_VDD_XI10.X0_PGD 6.1888e-19
cc_5 N_VSS_XI7.X0_S N_VDD_XI8.X0_S 4.21365e-19
cc_6 N_VSS_c_6_p N_VDD_XI8.X0_S 3.8999e-19
cc_7 N_VSS_XI8.X0_PGD N_VDD_XI7.X0_PGD 5.98857e-19
cc_8 N_VSS_c_8_p N_VDD_c_87_n 6.35797e-19
cc_9 N_VSS_c_9_p N_VDD_c_88_n 2.61781e-19
cc_10 N_VSS_c_10_p N_VDD_c_88_n 0.00161042f
cc_11 N_VSS_c_11_p N_VDD_c_88_n 0.00118088f
cc_12 N_VSS_c_12_p N_VDD_c_88_n 0.00296683f
cc_13 N_VSS_c_13_p N_VDD_c_88_n 0.00183744f
cc_14 N_VSS_c_9_p N_VDD_c_93_n 9.27292e-19
cc_15 N_VSS_c_15_p N_VDD_c_93_n 3.72495e-19
cc_16 N_VSS_c_16_p N_VDD_c_93_n 8.87931e-19
cc_17 N_VSS_c_10_p N_VDD_c_93_n 9.0356e-19
cc_18 N_VSS_c_11_p N_VDD_c_93_n 4.3265e-19
cc_19 N_VSS_c_19_p N_VDD_c_93_n 3.0156e-19
cc_20 N_VSS_c_12_p N_VDD_c_99_n 0.00167687f
cc_21 N_VSS_c_10_p N_VDD_c_100_n 0.00121886f
cc_22 N_VSS_c_19_p N_VDD_c_100_n 3.71304e-19
cc_23 N_VSS_XI6.X0_S N_VDD_c_102_n 4.24828e-19
cc_24 N_VSS_c_24_p N_VDD_c_102_n 0.00115189f
cc_25 N_VSS_c_2_p N_VDD_c_102_n 4.59126e-19
cc_26 N_VSS_c_24_p N_VDD_c_105_n 9.72233e-19
cc_27 N_VSS_c_27_p N_VDD_c_105_n 8.14547e-19
cc_28 N_VSS_c_28_p N_VDD_c_105_n 3.32851e-19
cc_29 N_VSS_XI7.X0_S N_VDD_c_108_n 3.8999e-19
cc_30 N_VSS_c_6_p N_VDD_c_108_n 5.78716e-19
cc_31 N_VSS_c_31_p N_VDD_c_108_n 0.00180659f
cc_32 N_VSS_c_10_p N_VDD_c_111_n 3.8999e-19
cc_33 N_VSS_c_11_p N_VDD_c_111_n 0.00181085f
cc_34 N_VSS_c_10_p N_Z_XI9.X0_D 8.835e-19
cc_35 N_VSS_c_11_p N_Z_XI9.X0_D 0.00246958f
cc_36 N_VSS_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_37 N_VSS_c_2_p N_Z_XI6.X0_D 3.48267e-19
cc_38 N_VSS_XI6.X0_S N_Z_XI10.X0_D 3.43419e-19
cc_39 N_VSS_XI7.X0_S N_Z_XI10.X0_D 3.43419e-19
cc_40 N_VSS_c_2_p N_Z_XI10.X0_D 3.48267e-19
cc_41 N_VSS_c_6_p N_Z_XI10.X0_D 3.48267e-19
cc_42 N_VSS_XI6.X0_S N_Z_c_170_n 3.48267e-19
cc_43 N_VSS_c_10_p N_Z_c_170_n 0.00217565f
cc_44 N_VSS_c_2_p N_Z_c_170_n 5.69026e-19
cc_45 N_VSS_c_11_p N_Z_c_170_n 8.835e-19
cc_46 N_VSS_c_12_p N_Z_c_170_n 7.10715e-19
cc_47 N_VSS_c_19_p N_Z_c_170_n 3.30259e-19
cc_48 N_VSS_XI6.X0_S N_Z_c_176_n 3.48267e-19
cc_49 N_VSS_XI7.X0_S N_Z_c_176_n 3.48267e-19
cc_50 N_VSS_c_2_p N_Z_c_176_n 5.69026e-19
cc_51 N_VSS_c_6_p N_Z_c_176_n 5.69026e-19
cc_52 N_VSS_c_2_p N_Z_c_180_n 0.00191849f
cc_53 N_VSS_c_12_p N_Z_c_180_n 5.57576e-19
cc_54 N_VSS_c_19_p N_Z_c_180_n 0.00201399f
cc_55 N_VSS_c_28_p N_Z_c_180_n 5.26184e-19
cc_56 N_VSS_XI9.X0_PGD N_C_c_212_n 4.30517e-19
cc_57 N_VSS_XI8.X0_PGD N_C_c_213_n 5.02359e-19
cc_58 N_VSS_c_28_p N_C_c_214_n 2.73385e-19
cc_59 N_VSS_XI9.X0_PGD N_C_c_215_n 4.3583e-19
cc_60 N_VSS_XI8.X0_PGD N_C_c_216_n 3.76133e-19
cc_61 N_VSS_c_61_p N_C_c_216_n 2.17009e-19
cc_62 N_VSS_XI9.X0_PGD N_B_XI9.X0_PGS 0.00109504f
cc_63 N_VSS_XI11.X0_PGD N_B_XI9.X0_PGS 2.15671e-19
cc_64 N_VSS_XI11.X0_PGD N_B_XI11.X0_PGS 0.00177732f
cc_65 N_VSS_XI8.X0_PGD N_B_XI11.X0_PGS 2.22194e-19
cc_66 N_VSS_c_61_p N_B_c_247_n 0.00177732f
cc_67 N_VSS_c_24_p N_B_c_248_n 0.00731987f
cc_68 N_VSS_c_16_p N_B_c_248_n 0.00109504f
cc_69 N_VSS_c_2_p B 2.11465e-19
cc_70 N_VSS_c_12_p B 2.74582e-19
cc_71 N_VSS_c_19_p B 2.99651e-19
cc_72 N_VSS_c_24_p N_A_XI11.X0_CG 2.66861e-19
cc_73 N_VSS_c_2_p N_A_c_272_n 3.13396e-19
cc_74 N_VSS_c_28_p N_A_c_272_n 5.88825e-19
cc_75 N_VSS_c_28_p A 5.88825e-19
cc_76 N_VSS_c_76_p A 2.39495e-19
cc_77 N_VSS_c_2_p N_A_c_276_n 0.00159849f
cc_78 N_VSS_c_28_p N_A_c_276_n 0.00924443f
cc_79 N_VSS_c_76_p N_A_c_276_n 5.12768e-19
cc_80 N_VDD_XI9.X0_S N_Z_XI9.X0_D 3.43419e-19
cc_81 N_VDD_c_93_n N_Z_XI9.X0_D 4.3265e-19
cc_82 N_VDD_c_102_n N_Z_XI9.X0_D 3.48267e-19
cc_83 N_VDD_c_100_n N_Z_XI6.X0_D 9.44213e-19
cc_84 N_VDD_c_111_n N_Z_XI6.X0_D 0.00246958f
cc_85 N_VDD_XI9.X0_S N_Z_XI11.X0_D 3.43419e-19
cc_86 N_VDD_XI8.X0_S N_Z_XI11.X0_D 3.43419e-19
cc_87 N_VDD_c_102_n N_Z_XI11.X0_D 3.48267e-19
cc_88 N_VDD_c_105_n N_Z_XI11.X0_D 4.3265e-19
cc_89 N_VDD_c_108_n N_Z_XI11.X0_D 3.72199e-19
cc_90 N_VDD_XI9.X0_S N_Z_c_170_n 3.48267e-19
cc_91 N_VDD_c_88_n N_Z_c_170_n 0.0013145f
cc_92 N_VDD_c_93_n N_Z_c_170_n 7.37531e-19
cc_93 N_VDD_c_100_n N_Z_c_170_n 0.00186578f
cc_94 N_VDD_c_102_n N_Z_c_170_n 7.73813e-19
cc_95 N_VDD_c_111_n N_Z_c_170_n 8.835e-19
cc_96 N_VDD_XI9.X0_S N_Z_c_176_n 3.48267e-19
cc_97 N_VDD_XI8.X0_S N_Z_c_176_n 3.48267e-19
cc_98 N_VDD_c_102_n N_Z_c_176_n 8.00908e-19
cc_99 N_VDD_c_105_n N_Z_c_176_n 5.78499e-19
cc_100 N_VDD_c_108_n N_Z_c_176_n 8.53368e-19
cc_101 N_VDD_c_93_n N_Z_c_180_n 8.36802e-19
cc_102 N_VDD_c_88_n C 2.63478e-19
cc_103 N_VDD_c_93_n C 0.00145322f
cc_104 N_VDD_c_102_n C 0.00155931f
cc_105 N_VDD_c_88_n N_C_c_214_n 2.14517e-19
cc_106 N_VDD_c_93_n N_C_c_214_n 8.61717e-19
cc_107 N_VDD_c_102_n N_C_c_214_n 0.00183615f
cc_108 N_VDD_c_105_n N_C_c_214_n 0.00557625f
cc_109 N_VDD_c_142_p N_C_c_214_n 5.42852e-19
cc_110 N_VDD_c_93_n N_C_c_215_n 7.51813e-19
cc_111 N_VDD_c_102_n N_C_c_215_n 8.66889e-19
cc_112 N_VDD_c_102_n N_C_c_216_n 2.22969e-19
cc_113 N_VDD_c_105_n N_C_c_216_n 2.63125e-19
cc_114 N_VDD_c_142_p N_C_c_216_n 3.66936e-19
cc_115 N_VDD_XI6.X0_PGD N_B_XI9.X0_PGS 0.00135245f
cc_116 N_VDD_XI10.X0_PGD N_B_XI9.X0_PGS 4.12959e-19
cc_117 N_VDD_c_150_p N_B_XI11.X0_PGS 0.00109105f
cc_118 N_VDD_c_150_p N_B_c_256_n 0.00258419f
cc_119 N_VDD_c_152_p N_B_c_256_n 4.12959e-19
cc_120 N_VDD_c_153_p N_B_c_258_n 0.00495207f
cc_121 N_VDD_c_111_n N_B_c_258_n 4.60491e-19
cc_122 N_VDD_XI10.X0_PGD N_A_XI11.X0_CG 4.83278e-19
cc_123 N_VDD_XI7.X0_PGD N_A_XI8.X0_PGS 0.00141985f
cc_124 N_VDD_c_105_n N_A_XI8.X0_PGS 2.26738e-19
cc_125 N_VDD_XI10.X0_PGD N_A_c_282_n 5.50272e-19
cc_126 N_VDD_XI7.X0_PGD N_A_c_283_n 3.23173e-19
cc_127 N_VDD_c_160_p N_A_c_283_n 0.00145458f
cc_128 N_VDD_c_152_p N_A_c_283_n 2.17009e-19
cc_129 N_Z_c_170_n N_C_c_212_n 6.18749e-19
cc_130 N_Z_c_176_n N_C_c_213_n 8.38264e-19
cc_131 N_Z_c_180_n N_C_c_214_n 0.0071108f
cc_132 N_Z_c_176_n N_A_XI11.X0_CG 2.49716e-19
cc_133 N_Z_c_176_n N_A_c_276_n 3.55289e-19
cc_134 N_Z_c_180_n N_A_c_276_n 0.00276659f
cc_135 N_C_c_212_n N_B_XI9.X0_PGS 0.00830899f
cc_136 N_C_c_215_n N_B_XI9.X0_PGS 3.76133e-19
cc_137 N_C_c_212_n N_B_XI11.X0_PGS 8.90713e-19
cc_138 N_C_c_213_n N_B_XI11.X0_PGS 5.42381e-19
cc_139 N_C_c_215_n N_B_c_258_n 3.15193e-19
cc_140 N_C_c_213_n N_A_XI11.X0_CG 0.0020589f
cc_141 N_C_c_213_n N_A_XI8.X0_PGS 0.00810452f
cc_142 N_C_c_214_n N_A_c_276_n 0.00121525f
cc_143 N_C_c_216_n N_A_c_283_n 3.16599e-19
cc_144 N_B_XI9.X0_PGS N_A_XI11.X0_CG 0.00106357f
cc_145 N_B_XI11.X0_PGS N_A_XI11.X0_CG 0.00765248f
cc_146 B N_A_c_272_n 3.39698e-19
cc_147 N_B_c_258_n N_A_c_272_n 3.48267e-19
cc_148 B N_A_c_282_n 3.48267e-19
cc_149 N_B_c_258_n N_A_c_282_n 5.15124e-19
*
.ends
*
*
.subckt MIN3_HPNW1 A B C Y VDD VSS
xgate (VSS VDD Y C B A) G3_MIN3_T6_N1
.ends
*
* File: G4_MUX2_N1.pex.netlist
* Created: Wed Mar  9 17:10:36 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MUX2_N1_VDD 2 4 6 8 10 12 14 18 20 38 49 58 84 85 87 89 93 95 96
+ 99 101 105 107 111 113 115 120 122 124 125 126 127 128 134 139 148 Vss
c140 148 Vss 0.00577129f
c141 139 Vss 0.00441689f
c142 134 Vss 0.00586273f
c143 128 Vss 3.56526e-19
c144 127 Vss 2.39889e-19
c145 126 Vss 4.22747e-19
c146 125 Vss 2.39889e-19
c147 122 Vss 0.00188211f
c148 120 Vss 0.00629792f
c149 115 Vss 0.00178287f
c150 113 Vss 0.00614865f
c151 111 Vss 6.94069e-19
c152 107 Vss 0.00775764f
c153 105 Vss 0.001258f
c154 101 Vss 0.00169538f
c155 99 Vss 4.33371e-19
c156 96 Vss 6.1175e-19
c157 95 Vss 0.00337348f
c158 93 Vss 0.00135966f
c159 89 Vss 0.00148319f
c160 87 Vss 0.00118366f
c161 85 Vss 0.00653402f
c162 84 Vss 0.00317212f
c163 83 Vss 0.00175227f
c164 59 Vss 0.0798032f
c165 58 Vss 0.102888f
c166 49 Vss 0.0346129f
c167 48 Vss 0.100303f
c168 39 Vss 0.0355046f
c169 38 Vss 0.100457f
c170 20 Vss 0.00271849f
c171 18 Vss 0.0807095f
c172 14 Vss 0.0816769f
c173 12 Vss 0.00155055f
c174 10 Vss 0.0815741f
c175 8 Vss 0.0807057f
c176 6 Vss 0.0842982f
c177 4 Vss 0.0825471f
c178 2 Vss 0.00231862f
r179 121 128 0.551426
r180 121 122 4.16786
r181 120 128 0.551426
r182 119 120 13.3371
r183 115 128 0.0828784
r184 115 117 1.82344
r185 114 127 0.494161
r186 113 119 0.652036
r187 113 114 10.1279
r188 111 148 1.16709
r189 109 127 0.128424
r190 109 111 2.16729
r191 108 126 0.494161
r192 107 122 0.652036
r193 107 108 13.0037
r194 103 126 0.128424
r195 103 105 4.83471
r196 102 125 0.494161
r197 101 127 0.494161
r198 101 102 4.58464
r199 99 139 1.16709
r200 97 125 0.128424
r201 97 99 2.16729
r202 95 126 0.494161
r203 95 96 7.46046
r204 93 134 1.16709
r205 91 96 0.652036
r206 91 93 2.16729
r207 87 89 1.82344
r208 86 124 0.326018
r209 85 125 0.494161
r210 85 86 10.1279
r211 84 87 0.655813
r212 83 124 0.326018
r213 83 84 4.16786
r214 64 148 0.238214
r215 64 66 1.92555
r216 59 66 0.5835
r217 58 60 0.652036
r218 58 59 2.8008
r219 55 66 0.0685365
r220 51 139 0.238214
r221 49 51 1.45875
r222 48 52 0.652036
r223 48 51 1.45875
r224 45 49 0.652036
r225 41 134 0.238214
r226 39 41 1.45875
r227 38 42 0.652036
r228 38 41 1.45875
r229 35 39 0.652036
r230 20 117 1.16709
r231 18 60 2.5674
r232 14 55 2.5674
r233 12 105 1.16709
r234 10 52 2.5674
r235 8 45 2.5674
r236 6 35 2.5674
r237 4 42 2.5674
r238 2 89 1.16709
.ends

.subckt PM_G4_MUX2_N1_VSS 2 4 6 8 10 12 16 18 20 38 39 48 49 51 59 84 89 94 99
+ 104 109 118 123 132 141 142 146 152 153 158 164 170 172 177 179 181 182 183
+ 184 185 Vss
c132 185 Vss 4.28045e-19
c133 184 Vss 3.62111e-19
c134 183 Vss 3.87529e-19
c135 182 Vss 3.75522e-19
c136 179 Vss 0.00396469f
c137 177 Vss 0.00140343f
c138 172 Vss 0.00128299f
c139 170 Vss 0.00250671f
c140 164 Vss 0.00572414f
c141 158 Vss 0.00417852f
c142 153 Vss 5.94991e-19
c143 152 Vss 0.00253786f
c144 146 Vss 0.00510722f
c145 142 Vss 0.00100335f
c146 141 Vss 0.00361314f
c147 132 Vss 0.00636077f
c148 123 Vss 0.00367258f
c149 118 Vss 0.0040616f
c150 109 Vss 3.31973e-19
c151 104 Vss 0.00116949f
c152 99 Vss 0.00135225f
c153 94 Vss 3.56537e-19
c154 89 Vss 8.02281e-19
c155 84 Vss 0.00135359f
c156 65 Vss 0.0785271f
c157 59 Vss 0.0340359f
c158 58 Vss 0.0688517f
c159 49 Vss 0.0338093f
c160 48 Vss 0.0993447f
c161 39 Vss 0.0341976f
c162 38 Vss 0.0984533f
c163 20 Vss 0.0819076f
c164 18 Vss 0.00227065f
c165 16 Vss 0.0807095f
c166 12 Vss 0.0827078f
c167 10 Vss 0.0826808f
c168 8 Vss 0.00150258f
c169 6 Vss 0.00290641f
c170 4 Vss 0.081612f
c171 2 Vss 0.0842992f
r172 178 185 0.551426
r173 178 179 13.3371
r174 177 185 0.551426
r175 176 177 4.16786
r176 172 185 0.0828784
r177 171 184 0.494161
r178 170 179 0.652036
r179 170 171 4.41793
r180 166 184 0.128424
r181 165 183 0.494161
r182 164 176 0.652036
r183 164 165 13.0037
r184 160 183 0.128424
r185 159 182 0.494161
r186 158 184 0.494161
r187 158 159 10.2946
r188 154 182 0.128424
r189 152 183 0.494161
r190 152 153 7.46046
r191 148 153 0.652036
r192 147 181 0.326018
r193 146 182 0.494161
r194 146 147 10.1279
r195 141 181 0.326018
r196 140 142 0.655813
r197 140 141 4.16786
r198 109 172 1.82344
r199 104 132 1.16709
r200 104 166 2.16729
r201 99 160 4.83471
r202 94 123 1.16709
r203 94 154 2.16729
r204 89 118 1.16709
r205 89 148 2.16729
r206 84 142 1.82344
r207 65 132 0.238214
r208 63 65 1.8672
r209 60 63 0.0685365
r210 58 63 0.5835
r211 58 59 2.8008
r212 55 59 0.652036
r213 51 123 0.238214
r214 49 51 1.45875
r215 48 52 0.652036
r216 48 51 1.45875
r217 45 49 0.652036
r218 41 118 0.238214
r219 39 41 1.45875
r220 38 42 0.652036
r221 38 41 1.45875
r222 35 39 0.652036
r223 20 60 2.5674
r224 18 109 1.16709
r225 16 55 2.5674
r226 12 52 2.5674
r227 10 45 2.5674
r228 8 99 1.16709
r229 6 84 1.16709
r230 4 42 2.5674
r231 2 35 2.5674
.ends

.subckt PM_G4_MUX2_N1_ZI 2 4 6 8 28 50 55 60 65 81 82 91 Vss
c67 82 Vss 9.74571e-19
c68 81 Vss 0.00289684f
c69 65 Vss 0.00556163f
c70 60 Vss 8.37584e-19
c71 55 Vss 0.00123466f
c72 50 Vss 0.00178991f
c73 28 Vss 0.206432f
c74 23 Vss 0.0247918f
c75 8 Vss 0.00143442f
c76 6 Vss 0.00143442f
c77 4 Vss 0.0815973f
c78 2 Vss 0.0715834f
r79 87 91 0.494161
r80 83 91 0.494161
r81 81 91 0.128424
r82 81 82 13.2121
r83 77 82 0.652036
r84 60 87 3.66771
r85 55 83 4.33457
r86 50 65 1.16709
r87 50 77 2.16729
r88 31 65 0.0476429
r89 29 31 0.326018
r90 29 31 0.1167
r91 28 32 0.652036
r92 28 31 6.7686
r93 27 65 0.357321
r94 23 31 0.326018
r95 23 27 0.40845
r96 8 60 1.16709
r97 6 55 1.16709
r98 4 32 2.5674
r99 2 27 2.15895
.ends

.subckt PM_G4_MUX2_N1_Z 2 18 Vss
c12 18 Vss 2.88294e-19
c13 2 Vss 0.00150258f
r14 2 18 1.16709
.ends

.subckt PM_G4_MUX2_N1_SELI 2 6 8 21 33 35 36 38 43 53 58 72 77 78 Vss
c81 78 Vss 6.39942e-19
c82 77 Vss 5.11483e-19
c83 72 Vss 0.00145166f
c84 58 Vss 0.0021541f
c85 53 Vss 0.00198421f
c86 43 Vss 9.80359e-19
c87 38 Vss 0.00153196f
c88 36 Vss 2.15854e-19
c89 35 Vss 0.00258645f
c90 33 Vss 0.00238155f
c91 21 Vss 0.0575125f
c92 6 Vss 0.0575499f
c93 2 Vss 0.00172036f
r94 77 78 0.655813
r95 76 77 3.501
r96 72 76 0.655813
r97 43 53 1.16709
r98 43 72 2.00578
r99 43 46 0.833571
r100 38 58 1.16709
r101 38 78 2.00578
r102 35 46 0.0685365
r103 35 36 7.46046
r104 31 36 0.652036
r105 31 33 5.58493
r106 21 58 0.50025
r107 18 53 0.50025
r108 8 21 1.80885
r109 6 18 1.80885
r110 2 33 1.16709
.ends

.subckt PM_G4_MUX2_N1_SEL 2 4 6 8 16 17 22 26 37 40 41 44 45 46 47 52 58 63 68
+ 73 Vss
c78 73 Vss 0.00176698f
c79 68 Vss 0.00182856f
c80 63 Vss 0.00250521f
c81 58 Vss 7.07944e-19
c82 52 Vss 2.9409e-19
c83 47 Vss 2.03369e-19
c84 46 Vss 3.54223e-19
c85 45 Vss 7.77909e-19
c86 44 Vss 0.00151239f
c87 41 Vss 0.00163463f
c88 37 Vss 0.00192905f
c89 26 Vss 0.0575125f
c90 22 Vss 0.0712295f
c91 20 Vss 0.0247918f
c92 17 Vss 0.0358042f
c93 16 Vss 0.175331f
c94 8 Vss 0.0575125f
c95 2 Vss 0.084915f
r96 58 73 1.16709
r97 58 60 0.5835
r98 55 68 1.16709
r99 52 55 0.5835
r100 50 63 1.16709
r101 47 50 0.5835
r102 45 60 0.0685365
r103 45 46 1.70882
r104 43 46 0.652036
r105 43 44 2.50071
r106 42 52 0.0685365
r107 41 44 0.652036
r108 41 42 1.70882
r109 38 47 0.0685365
r110 38 40 1.62546
r111 37 52 0.0685365
r112 37 40 2.95918
r113 36 63 0.0476429
r114 33 73 0.50025
r115 26 68 0.50025
r116 22 63 0.357321
r117 20 36 0.326018
r118 20 22 0.40845
r119 17 36 6.7686
r120 16 36 0.326018
r121 16 36 0.1167
r122 13 17 0.652036
r123 8 33 1.80885
r124 6 26 1.80885
r125 4 22 2.15895
r126 2 13 2.5674
.ends

.subckt PM_G4_MUX2_N1_B 2 4 14 20 23 Vss
c31 23 Vss 0.00482401f
c32 20 Vss 4.63929e-19
c33 14 Vss 0.0843809f
c34 2 Vss 0.446304f
r35 17 23 1.16709
r36 17 20 0.0364688
r37 14 23 0.238214
r38 11 14 1.92555
r39 7 11 0.0685365
r40 4 7 2.5674
r41 2 4 12.837
.ends

.subckt PM_G4_MUX2_N1_A 2 4 14 20 23 Vss
c25 23 Vss 0.00557714f
c26 20 Vss 2.81445e-19
c27 14 Vss 0.0830192f
c28 2 Vss 0.44929f
r29 17 23 1.16709
r30 17 20 0.0729375
r31 12 23 0.238214
r32 12 14 1.92555
r33 7 14 0.0685365
r34 2 4 12.837
r35 2 7 2.5674
.ends

.subckt G4_MUX2_N1  VDD VSS Z SEL B A
*
* A	A
* B	B
* SEL	SEL
* Z	Z
* VSS	VSS
* VDD	VDD
XI7.X0 N_VDD_XI7.X0_D N_VSS_XI7.X0_PGD N_ZI_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_Z_XI7.X0_S TIGFET_HPNW1
XI1.X0 N_SELI_XI1.X0_D N_VDD_XI1.X0_PGD N_SEL_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
XI6.X0 N_Z_XI7.X0_S N_VDD_XI6.X0_PGD N_ZI_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW1
XI2.X0 N_SELI_XI1.X0_D N_VSS_XI2.X0_PGD N_SEL_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI5.X0 N_ZI_XI5.X0_D N_VDD_XI5.X0_PGD N_SELI_XI5.X0_CG N_B_XI5.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW1
XI3.X0 N_ZI_XI3.X0_D N_VSS_XI3.X0_PGD N_SEL_XI3.X0_CG N_B_XI3.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI4.X0 N_ZI_XI5.X0_D N_VDD_XI4.X0_PGD N_SEL_XI4.X0_CG N_A_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW1
XI0.X0 N_ZI_XI3.X0_D N_VSS_XI0.X0_PGD N_SELI_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW1
*
x_PM_G4_MUX2_N1_VDD N_VDD_XI7.X0_D N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS
+ N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI2.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_14_p N_VDD_c_11_p N_VDD_c_136_p
+ N_VDD_c_18_p N_VDD_c_12_p N_VDD_c_46_p N_VDD_c_17_p N_VDD_c_22_p N_VDD_c_15_p
+ N_VDD_c_48_p N_VDD_c_20_p N_VDD_c_3_p N_VDD_c_6_p N_VDD_c_16_p N_VDD_c_28_p
+ N_VDD_c_8_p N_VDD_c_34_p N_VDD_c_9_p N_VDD_c_32_p VDD N_VDD_c_51_p
+ N_VDD_c_55_p N_VDD_c_58_p N_VDD_c_65_p N_VDD_c_25_p N_VDD_c_21_p N_VDD_c_95_p
+ Vss PM_G4_MUX2_N1_VDD
x_PM_G4_MUX2_N1_VSS N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS N_VSS_XI1.X0_S
+ N_VSS_XI6.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS N_VSS_XI3.X0_PGD
+ N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_151_n N_VSS_c_153_n N_VSS_c_265_p
+ N_VSS_c_154_n N_VSS_c_257_p N_VSS_c_156_n N_VSS_c_157_n N_VSS_c_158_n
+ N_VSS_c_162_n N_VSS_c_166_n N_VSS_c_170_n N_VSS_c_173_n N_VSS_c_176_n
+ N_VSS_c_180_n N_VSS_c_184_n N_VSS_c_185_n N_VSS_c_186_n N_VSS_c_187_n
+ N_VSS_c_189_n N_VSS_c_192_n N_VSS_c_193_n N_VSS_c_196_n N_VSS_c_199_n
+ N_VSS_c_200_n N_VSS_c_201_n N_VSS_c_202_n VSS N_VSS_c_206_n N_VSS_c_207_n
+ N_VSS_c_208_n N_VSS_c_209_n Vss PM_G4_MUX2_N1_VSS
x_PM_G4_MUX2_N1_ZI N_ZI_XI7.X0_CG N_ZI_XI6.X0_CG N_ZI_XI5.X0_D N_ZI_XI3.X0_D
+ N_ZI_c_278_n N_ZI_c_294_n N_ZI_c_280_n N_ZI_c_282_n N_ZI_c_287_n N_ZI_c_288_n
+ N_ZI_c_311_n N_ZI_c_326_p Vss PM_G4_MUX2_N1_ZI
x_PM_G4_MUX2_N1_Z N_Z_XI7.X0_S Z Vss PM_G4_MUX2_N1_Z
x_PM_G4_MUX2_N1_SELI N_SELI_XI1.X0_D N_SELI_XI5.X0_CG N_SELI_XI0.X0_CG
+ N_SELI_c_371_n N_SELI_c_356_n N_SELI_c_359_n N_SELI_c_387_n N_SELI_c_364_n
+ N_SELI_c_365_n N_SELI_c_367_n N_SELI_c_379_n N_SELI_c_381_n N_SELI_c_395_n
+ N_SELI_c_398_n Vss PM_G4_MUX2_N1_SELI
x_PM_G4_MUX2_N1_SEL N_SEL_XI1.X0_CG N_SEL_XI2.X0_CG N_SEL_XI3.X0_CG
+ N_SEL_XI4.X0_CG N_SEL_c_434_n N_SEL_c_460_n N_SEL_c_449_n N_SEL_c_495_p
+ N_SEL_c_436_n SEL N_SEL_c_438_n N_SEL_c_439_n N_SEL_c_440_n N_SEL_c_465_n
+ N_SEL_c_453_n N_SEL_c_468_n N_SEL_c_442_n N_SEL_c_443_n N_SEL_c_444_n
+ N_SEL_c_445_n Vss PM_G4_MUX2_N1_SEL
x_PM_G4_MUX2_N1_B N_B_XI5.X0_PGS N_B_XI3.X0_PGS N_B_c_518_n B N_B_c_514_n Vss
+ PM_G4_MUX2_N1_B
x_PM_G4_MUX2_N1_A N_A_XI4.X0_PGS N_A_XI0.X0_PGS N_A_c_544_n A N_A_c_550_n Vss
+ PM_G4_MUX2_N1_A
cc_1 N_VDD_XI1.X0_PGS N_VSS_XI7.X0_PGD 2.27468e-19
cc_2 N_VDD_XI6.X0_PGD N_VSS_XI7.X0_PGS 0.00173038f
cc_3 N_VDD_c_3_p N_VSS_XI6.X0_S 3.7884e-19
cc_4 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.0016786f
cc_5 N_VDD_XI6.X0_PGS N_VSS_XI2.X0_PGS 2.11937e-19
cc_6 N_VDD_c_6_p N_VSS_XI2.X0_PGS 2.56778e-19
cc_7 N_VDD_XI5.X0_PGD N_VSS_XI3.X0_PGD 2.1536e-19
cc_8 N_VDD_c_8_p N_VSS_XI4.X0_S 3.7884e-19
cc_9 N_VDD_c_9_p N_VSS_XI4.X0_S 9.5668e-19
cc_10 N_VDD_XI4.X0_PGD N_VSS_XI0.X0_PGD 2.1536e-19
cc_11 N_VDD_c_11_p N_VSS_c_151_n 0.00173038f
cc_12 N_VDD_c_12_p N_VSS_c_151_n 3.60588e-19
cc_13 N_VDD_c_12_p N_VSS_c_153_n 3.80388e-19
cc_14 N_VDD_c_14_p N_VSS_c_154_n 0.0016786f
cc_15 N_VDD_c_15_p N_VSS_c_154_n 2.72324e-19
cc_16 N_VDD_c_16_p N_VSS_c_156_n 8.01165e-19
cc_17 N_VDD_c_17_p N_VSS_c_157_n 9.30123e-19
cc_18 N_VDD_c_18_p N_VSS_c_158_n 8.69498e-19
cc_19 N_VDD_c_12_p N_VSS_c_158_n 0.00141228f
cc_20 N_VDD_c_20_p N_VSS_c_158_n 8.51944e-19
cc_21 N_VDD_c_21_p N_VSS_c_158_n 3.48267e-19
cc_22 N_VDD_c_22_p N_VSS_c_162_n 8.56577e-19
cc_23 N_VDD_c_15_p N_VSS_c_162_n 0.00141228f
cc_24 N_VDD_c_6_p N_VSS_c_162_n 0.00181129f
cc_25 N_VDD_c_25_p N_VSS_c_162_n 3.48267e-19
cc_26 N_VDD_c_20_p N_VSS_c_166_n 3.92901e-19
cc_27 N_VDD_c_3_p N_VSS_c_166_n 4.58491e-19
cc_28 N_VDD_c_28_p N_VSS_c_166_n 7.06793e-19
cc_29 N_VDD_c_9_p N_VSS_c_166_n 2.71563e-19
cc_30 N_VDD_c_6_p N_VSS_c_170_n 2.93442e-19
cc_31 N_VDD_c_16_p N_VSS_c_170_n 0.00161703f
cc_32 N_VDD_c_32_p N_VSS_c_170_n 4.6996e-19
cc_33 N_VDD_c_8_p N_VSS_c_173_n 4.73473e-19
cc_34 N_VDD_c_34_p N_VSS_c_173_n 2.13058e-19
cc_35 N_VDD_c_9_p N_VSS_c_173_n 0.00165395f
cc_36 N_VDD_c_18_p N_VSS_c_176_n 3.66936e-19
cc_37 N_VDD_c_12_p N_VSS_c_176_n 0.00112249f
cc_38 N_VDD_c_20_p N_VSS_c_176_n 3.99794e-19
cc_39 N_VDD_c_21_p N_VSS_c_176_n 8.07896e-19
cc_40 N_VDD_c_22_p N_VSS_c_180_n 3.82294e-19
cc_41 N_VDD_c_15_p N_VSS_c_180_n 0.00112249f
cc_42 N_VDD_c_6_p N_VSS_c_180_n 9.55349e-19
cc_43 N_VDD_c_25_p N_VSS_c_180_n 8.0279e-19
cc_44 N_VDD_c_16_p N_VSS_c_184_n 2.03837e-19
cc_45 N_VDD_c_22_p N_VSS_c_185_n 3.85245e-19
cc_46 N_VDD_c_46_p N_VSS_c_186_n 4.93614e-19
cc_47 N_VDD_c_15_p N_VSS_c_187_n 0.003995f
cc_48 N_VDD_c_48_p N_VSS_c_187_n 0.00163298f
cc_49 N_VDD_c_12_p N_VSS_c_189_n 0.00401122f
cc_50 N_VDD_c_3_p N_VSS_c_189_n 0.0013091f
cc_51 N_VDD_c_51_p N_VSS_c_189_n 0.0010079f
cc_52 N_VDD_c_12_p N_VSS_c_192_n 0.00176255f
cc_53 N_VDD_c_15_p N_VSS_c_193_n 0.00131941f
cc_54 N_VDD_c_16_p N_VSS_c_193_n 0.00593836f
cc_55 N_VDD_c_55_p N_VSS_c_193_n 0.00111239f
cc_56 N_VDD_c_3_p N_VSS_c_196_n 0.0013091f
cc_57 N_VDD_c_8_p N_VSS_c_196_n 0.00841532f
cc_58 N_VDD_c_58_p N_VSS_c_196_n 9.6871e-19
cc_59 N_VDD_c_16_p N_VSS_c_199_n 0.00454933f
cc_60 N_VDD_c_34_p N_VSS_c_200_n 5.34009e-19
cc_61 N_VDD_c_9_p N_VSS_c_201_n 0.00304617f
cc_62 N_VDD_c_6_p N_VSS_c_202_n 2.5062e-19
cc_63 N_VDD_c_9_p N_VSS_c_202_n 0.00529507f
cc_64 N_VDD_c_32_p N_VSS_c_202_n 0.00267625f
cc_65 N_VDD_c_65_p N_VSS_c_202_n 0.0010706f
cc_66 N_VDD_c_15_p N_VSS_c_206_n 7.74609e-19
cc_67 N_VDD_c_3_p N_VSS_c_207_n 0.00104966f
cc_68 N_VDD_c_16_p N_VSS_c_208_n 7.61747e-19
cc_69 N_VDD_c_9_p N_VSS_c_209_n 8.91588e-19
cc_70 N_VDD_c_21_p N_ZI_XI6.X0_CG 9.92565e-19
cc_71 N_VDD_XI2.X0_S N_ZI_XI3.X0_D 3.43419e-19
cc_72 N_VDD_XI0.X0_S N_ZI_XI3.X0_D 3.43419e-19
cc_73 N_VDD_c_6_p N_ZI_XI3.X0_D 3.48267e-19
cc_74 N_VDD_c_34_p N_ZI_XI3.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_PGD N_ZI_c_278_n 2.22031e-19
cc_76 N_VDD_XI6.X0_PGD N_ZI_c_278_n 3.91104e-19
cc_77 N_VDD_c_8_p N_ZI_c_280_n 5.01863e-19
cc_78 N_VDD_c_9_p N_ZI_c_280_n 4.66891e-19
cc_79 N_VDD_XI2.X0_S N_ZI_c_282_n 3.48267e-19
cc_80 N_VDD_XI0.X0_S N_ZI_c_282_n 3.48267e-19
cc_81 N_VDD_c_6_p N_ZI_c_282_n 4.97272e-19
cc_82 N_VDD_c_16_p N_ZI_c_282_n 5.01863e-19
cc_83 N_VDD_c_34_p N_ZI_c_282_n 5.226e-19
cc_84 N_VDD_c_25_p N_ZI_c_287_n 5.3845e-19
cc_85 N_VDD_c_15_p N_ZI_c_288_n 3.65425e-19
cc_86 N_VDD_XI7.X0_D N_Z_XI7.X0_S 3.43419e-19
cc_87 N_VDD_c_12_p N_Z_XI7.X0_S 3.7884e-19
cc_88 N_VDD_c_17_p N_Z_XI7.X0_S 3.72199e-19
cc_89 N_VDD_XI7.X0_D Z 3.48267e-19
cc_90 N_VDD_c_12_p Z 5.12447e-19
cc_91 N_VDD_c_17_p Z 7.4527e-19
cc_92 N_VDD_XI2.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_93 N_VDD_c_15_p N_SELI_XI1.X0_D 3.7884e-19
cc_94 N_VDD_c_6_p N_SELI_XI1.X0_D 3.48267e-19
cc_95 N_VDD_c_95_p N_SELI_XI5.X0_CG 0.00237871f
cc_96 N_VDD_XI2.X0_S N_SELI_c_356_n 3.48267e-19
cc_97 N_VDD_c_15_p N_SELI_c_356_n 5.34458e-19
cc_98 N_VDD_c_6_p N_SELI_c_356_n 6.883e-19
cc_99 N_VDD_XI6.X0_PGD N_SELI_c_359_n 2.27908e-19
cc_100 N_VDD_c_15_p N_SELI_c_359_n 2.61043e-19
cc_101 N_VDD_c_20_p N_SELI_c_359_n 5.3241e-19
cc_102 N_VDD_c_3_p N_SELI_c_359_n 2.36369e-19
cc_103 N_VDD_c_21_p N_SELI_c_359_n 3.99122e-19
cc_104 N_VDD_c_9_p N_SELI_c_364_n 4.30008e-19
cc_105 N_VDD_c_28_p N_SELI_c_365_n 7.54639e-19
cc_106 N_VDD_c_95_p N_SELI_c_365_n 5.0614e-19
cc_107 N_VDD_c_28_p N_SELI_c_367_n 4.85469e-19
cc_108 N_VDD_c_95_p N_SELI_c_367_n 0.0014909f
cc_109 N_VDD_c_25_p N_SEL_XI1.X0_CG 9.92565e-19
cc_110 N_VDD_XI1.X0_PGD N_SEL_c_434_n 4.04053e-19
cc_111 N_VDD_XI6.X0_PGD N_SEL_c_434_n 2.07349e-19
cc_112 N_VDD_XI2.X0_S N_SEL_c_436_n 9.18655e-19
cc_113 N_VDD_c_6_p N_SEL_c_436_n 0.00151457f
cc_114 N_VDD_c_16_p N_SEL_c_438_n 4.35337e-19
cc_115 N_VDD_c_9_p N_SEL_c_439_n 4.25334e-19
cc_116 N_VDD_c_16_p N_SEL_c_440_n 2.49768e-19
cc_117 N_VDD_c_8_p N_SEL_c_440_n 4.35337e-19
cc_118 N_VDD_c_9_p N_SEL_c_442_n 8.17234e-19
cc_119 N_VDD_c_21_p N_SEL_c_443_n 4.93609e-19
cc_120 N_VDD_c_95_p N_SEL_c_444_n 2.00604e-19
cc_121 N_VDD_XI4.X0_PGD N_SEL_c_445_n 3.11814e-19
cc_122 N_VDD_c_9_p N_SEL_c_445_n 3.66936e-19
cc_123 N_VDD_c_6_p N_B_XI5.X0_PGS 2.48132e-19
cc_124 N_VDD_c_6_p B 0.0014278f
cc_125 N_VDD_c_16_p B 0.00141439f
cc_126 N_VDD_c_6_p N_B_c_514_n 9.67317e-19
cc_127 N_VDD_c_16_p N_B_c_514_n 0.00117371f
cc_128 N_VDD_XI4.X0_PGD N_A_XI4.X0_PGS 0.00162178f
cc_129 N_VDD_c_9_p N_A_XI4.X0_PGS 9.35727e-19
cc_130 N_VDD_c_8_p N_A_c_544_n 3.3974e-19
cc_131 N_VDD_c_9_p N_A_c_544_n 4.15738e-19
cc_132 N_VDD_c_28_p A 5.43314e-19
cc_133 N_VDD_c_8_p A 0.00141439f
cc_134 N_VDD_c_9_p A 5.30212e-19
cc_135 N_VDD_c_95_p A 3.48267e-19
cc_136 N_VDD_c_136_p N_A_c_550_n 0.00480616f
cc_137 N_VDD_c_28_p N_A_c_550_n 4.04186e-19
cc_138 N_VDD_c_8_p N_A_c_550_n 0.00117371f
cc_139 N_VDD_c_9_p N_A_c_550_n 3.66936e-19
cc_140 N_VDD_c_95_p N_A_c_550_n 6.39485e-19
cc_141 N_VSS_c_176_n N_ZI_XI7.X0_CG 0.00234241f
cc_142 N_VSS_XI6.X0_S N_ZI_XI5.X0_D 3.43419e-19
cc_143 N_VSS_XI4.X0_S N_ZI_XI5.X0_D 3.43419e-19
cc_144 N_VSS_c_173_n N_ZI_XI5.X0_D 3.48267e-19
cc_145 N_VSS_XI7.X0_PGS N_ZI_c_278_n 3.99472e-19
cc_146 N_VSS_c_158_n N_ZI_c_294_n 0.00126951f
cc_147 N_VSS_c_176_n N_ZI_c_294_n 8.72558e-19
cc_148 N_VSS_XI6.X0_S N_ZI_c_280_n 3.48267e-19
cc_149 N_VSS_XI4.X0_S N_ZI_c_280_n 3.48267e-19
cc_150 N_VSS_c_166_n N_ZI_c_280_n 0.00100597f
cc_151 N_VSS_c_173_n N_ZI_c_280_n 4.40384e-19
cc_152 N_VSS_c_196_n N_ZI_c_280_n 5.12922e-19
cc_153 N_VSS_c_200_n N_ZI_c_280_n 6.1924e-19
cc_154 N_VSS_c_202_n N_ZI_c_280_n 0.00113121f
cc_155 N_VSS_c_193_n N_ZI_c_282_n 5.12922e-19
cc_156 N_VSS_c_158_n N_ZI_c_287_n 4.56568e-19
cc_157 N_VSS_c_176_n N_ZI_c_287_n 0.0014909f
cc_158 N_VSS_c_162_n N_ZI_c_288_n 4.17431e-19
cc_159 N_VSS_c_166_n N_ZI_c_288_n 6.40656e-19
cc_160 N_VSS_c_189_n N_ZI_c_288_n 0.00101727f
cc_161 N_VSS_c_193_n N_ZI_c_288_n 0.00147997f
cc_162 N_VSS_c_196_n N_ZI_c_288_n 2.59546e-19
cc_163 N_VSS_c_187_n N_ZI_c_311_n 0.0011789f
cc_164 N_VSS_XI6.X0_S N_Z_XI7.X0_S 3.43419e-19
cc_165 N_VSS_c_166_n N_Z_XI7.X0_S 3.48267e-19
cc_166 N_VSS_XI6.X0_S Z 3.48267e-19
cc_167 N_VSS_c_166_n Z 7.85754e-19
cc_168 N_VSS_XI1.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_169 N_VSS_c_157_n N_SELI_XI1.X0_D 3.48267e-19
cc_170 N_VSS_c_184_n N_SELI_c_371_n 0.00234241f
cc_171 N_VSS_c_157_n N_SELI_c_356_n 6.0686e-19
cc_172 N_VSS_c_166_n N_SELI_c_359_n 0.00130595f
cc_173 N_VSS_c_189_n N_SELI_c_359_n 4.10258e-19
cc_174 N_VSS_c_170_n N_SELI_c_364_n 0.00135778f
cc_175 N_VSS_c_184_n N_SELI_c_364_n 4.99367e-19
cc_176 N_VSS_c_196_n N_SELI_c_364_n 4.69529e-19
cc_177 N_VSS_c_202_n N_SELI_c_364_n 9.62347e-19
cc_178 N_VSS_c_170_n N_SELI_c_379_n 4.56568e-19
cc_179 N_VSS_c_184_n N_SELI_c_379_n 0.0014909f
cc_180 N_VSS_c_196_n N_SELI_c_381_n 7.6099e-19
cc_181 N_VSS_c_202_n N_SELI_c_381_n 6.2582e-19
cc_182 N_VSS_XI7.X0_PGS N_SEL_c_434_n 2.22031e-19
cc_183 N_VSS_XI2.X0_PGD N_SEL_c_434_n 3.91879e-19
cc_184 N_VSS_c_180_n N_SEL_c_449_n 0.00272336f
cc_185 N_VSS_c_193_n N_SEL_c_436_n 4.08267e-19
cc_186 N_VSS_c_202_n N_SEL_c_439_n 2.03139e-19
cc_187 N_VSS_c_196_n N_SEL_c_440_n 2.53418e-19
cc_188 N_VSS_c_257_p N_SEL_c_453_n 3.73191e-19
cc_189 N_VSS_c_162_n N_SEL_c_453_n 6.21258e-19
cc_190 N_VSS_c_162_n N_SEL_c_443_n 4.56568e-19
cc_191 N_VSS_c_180_n N_SEL_c_443_n 0.0014909f
cc_192 N_VSS_XI3.X0_PGD N_SEL_c_444_n 3.11814e-19
cc_193 N_VSS_c_184_n N_SEL_c_445_n 2.00604e-19
cc_194 N_VSS_XI2.X0_PGS N_B_XI5.X0_PGS 0.00172969f
cc_195 N_VSS_XI3.X0_PGD N_B_XI5.X0_PGS 0.00152606f
cc_196 N_VSS_c_265_p N_B_c_518_n 0.00172969f
cc_197 N_VSS_c_170_n B 3.98896e-19
cc_198 N_VSS_c_184_n B 3.5189e-19
cc_199 N_VSS_c_156_n N_B_c_514_n 0.00295829f
cc_200 N_VSS_c_170_n N_B_c_514_n 3.5189e-19
cc_201 N_VSS_c_180_n N_B_c_514_n 7.89771e-19
cc_202 N_VSS_c_184_n N_B_c_514_n 6.80896e-19
cc_203 N_VSS_c_196_n A 2.11858e-19
cc_204 N_ZI_c_282_n N_SELI_c_356_n 3.26181e-19
cc_205 N_ZI_c_288_n N_SELI_c_356_n 0.00213954f
cc_206 N_ZI_c_278_n N_SELI_c_359_n 4.92356e-19
cc_207 N_ZI_c_288_n N_SELI_c_359_n 0.00182433f
cc_208 N_ZI_c_278_n N_SELI_c_387_n 2.38253e-19
cc_209 N_ZI_c_294_n N_SELI_c_387_n 0.00150231f
cc_210 N_ZI_c_287_n N_SELI_c_387_n 0.00110082f
cc_211 N_ZI_c_282_n N_SELI_c_364_n 0.00173524f
cc_212 N_ZI_c_280_n N_SELI_c_365_n 0.00183505f
cc_213 N_ZI_c_288_n N_SELI_c_365_n 0.00144518f
cc_214 N_ZI_c_280_n N_SELI_c_381_n 7.38292e-19
cc_215 N_ZI_c_288_n N_SELI_c_381_n 7.7914e-19
cc_216 N_ZI_c_280_n N_SELI_c_395_n 5.82645e-19
cc_217 N_ZI_c_282_n N_SELI_c_395_n 3.22755e-19
cc_218 N_ZI_c_326_p N_SELI_c_395_n 6.45182e-19
cc_219 N_ZI_c_282_n N_SELI_c_398_n 7.64986e-19
cc_220 N_ZI_c_278_n N_SEL_c_434_n 0.00371647f
cc_221 N_ZI_c_287_n N_SEL_c_460_n 3.81736e-19
cc_222 N_ZI_XI3.X0_D N_SEL_c_438_n 9.94581e-19
cc_223 N_ZI_c_282_n N_SEL_c_438_n 0.00247421f
cc_224 N_ZI_c_280_n N_SEL_c_439_n 6.15647e-19
cc_225 N_ZI_c_326_p N_SEL_c_439_n 0.00107464f
cc_226 N_ZI_XI5.X0_D N_SEL_c_465_n 9.94581e-19
cc_227 N_ZI_c_280_n N_SEL_c_465_n 0.00243387f
cc_228 N_ZI_c_288_n N_SEL_c_453_n 0.00217047f
cc_229 N_ZI_c_282_n N_SEL_c_468_n 2.25033e-19
cc_230 N_ZI_c_278_n N_SEL_c_443_n 3.81736e-19
cc_231 N_ZI_XI6.X0_CG N_B_XI5.X0_PGS 0.00182649f
cc_232 N_Z_XI7.X0_S N_SELI_c_387_n 9.09799e-19
cc_233 Z N_SELI_c_387_n 0.00147087f
cc_234 N_SELI_c_356_n N_SEL_c_434_n 8.51271e-19
cc_235 N_SELI_c_365_n N_SEL_c_436_n 0.00269197f
cc_236 N_SELI_c_364_n N_SEL_c_438_n 0.00117605f
cc_237 N_SELI_c_356_n N_SEL_c_439_n 2.52418e-19
cc_238 N_SELI_c_364_n N_SEL_c_440_n 3.73414e-19
cc_239 N_SELI_c_365_n N_SEL_c_465_n 0.00160262f
cc_240 N_SELI_c_367_n N_SEL_c_465_n 9.78333e-19
cc_241 N_SELI_c_356_n N_SEL_c_453_n 0.00246582f
cc_242 N_SELI_c_359_n N_SEL_c_453_n 0.00269197f
cc_243 N_SELI_c_364_n N_SEL_c_468_n 2.32653e-19
cc_244 N_SELI_c_379_n N_SEL_c_468_n 3.48267e-19
cc_245 N_SELI_c_364_n N_SEL_c_442_n 9.4965e-19
cc_246 N_SELI_c_365_n N_SEL_c_442_n 2.32653e-19
cc_247 N_SELI_c_367_n N_SEL_c_442_n 3.48267e-19
cc_248 N_SELI_c_356_n N_SEL_c_443_n 9.71051e-19
cc_249 N_SELI_c_359_n N_SEL_c_443_n 6.26941e-19
cc_250 N_SELI_c_364_n N_SEL_c_444_n 3.48267e-19
cc_251 N_SELI_c_365_n N_SEL_c_444_n 7.22902e-19
cc_252 N_SELI_c_367_n N_SEL_c_444_n 0.0049864f
cc_253 N_SELI_c_379_n N_SEL_c_444_n 9.11855e-19
cc_254 N_SELI_c_364_n N_SEL_c_445_n 4.99367e-19
cc_255 N_SELI_c_365_n N_SEL_c_445_n 3.68647e-19
cc_256 N_SELI_c_367_n N_SEL_c_445_n 9.28301e-19
cc_257 N_SELI_c_379_n N_SEL_c_445_n 0.00490516f
cc_258 N_SELI_XI5.X0_CG N_B_XI5.X0_PGS 4.41254e-19
cc_259 N_SELI_c_356_n N_B_XI5.X0_PGS 2.21243e-19
cc_260 N_SELI_c_359_n N_B_XI5.X0_PGS 7.89402e-19
cc_261 N_SELI_c_367_n N_B_XI5.X0_PGS 0.00186882f
cc_262 N_SELI_c_367_n N_B_c_514_n 2.00604e-19
cc_263 N_SELI_c_371_n N_A_XI4.X0_PGS 4.65768e-19
cc_264 N_SELI_c_379_n N_A_XI4.X0_PGS 0.00276355f
cc_265 N_SELI_c_379_n N_A_c_550_n 2.00604e-19
cc_266 N_SEL_c_449_n N_B_XI5.X0_PGS 2.07014e-19
cc_267 N_SEL_c_495_p N_B_XI5.X0_PGS 4.3669e-19
cc_268 N_SEL_c_436_n N_B_XI5.X0_PGS 7.4877e-19
cc_269 N_SEL_c_443_n N_B_XI5.X0_PGS 0.00100354f
cc_270 N_SEL_c_444_n N_B_XI5.X0_PGS 0.00202689f
cc_271 N_SEL_c_468_n B 6.87706e-19
cc_272 N_SEL_c_444_n B 4.56568e-19
cc_273 N_SEL_c_495_p N_B_c_514_n 0.00234241f
cc_274 N_SEL_c_468_n N_B_c_514_n 5.02946e-19
cc_275 N_SEL_c_444_n N_B_c_514_n 0.0014909f
cc_276 N_SEL_XI4.X0_CG N_A_XI4.X0_PGS 4.54863e-19
cc_277 N_SEL_c_445_n N_A_XI4.X0_PGS 0.00276355f
cc_278 N_SEL_c_442_n A 7.05846e-19
cc_279 N_SEL_c_445_n A 4.56568e-19
cc_280 N_SEL_XI4.X0_CG N_A_c_550_n 0.00234241f
cc_281 N_SEL_c_442_n N_A_c_550_n 5.02946e-19
cc_282 N_SEL_c_445_n N_A_c_550_n 0.0014909f
cc_283 N_B_XI5.X0_PGS N_A_XI4.X0_PGS 0.00137635f
*
.ends
*
*
.subckt MUX2_HPNW1 A B S0 Y VDD VSS
xgate (VDD VSS Y S0 B A) G4_MUX2_N1
.ends
*
* File: G3_MUXI2_N1.pex.netlist
* Created: Wed Mar  9 13:36:32 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MUXI2_N1_VSS 2 4 6 8 10 12 14 29 31 39 63 68 73 78 83 92 101 110
+ 115 121 127 133 135 140 142 144 145 146 147 Vss
c86 147 Vss 4.28045e-19
c87 146 Vss 3.62111e-19
c88 145 Vss 3.75522e-19
c89 142 Vss 0.00430383f
c90 140 Vss 0.00143623f
c91 135 Vss 0.00139741f
c92 133 Vss 0.002505f
c93 128 Vss 0.00127887f
c94 127 Vss 0.00644124f
c95 121 Vss 0.00399642f
c96 116 Vss 0.0013489f
c97 115 Vss 0.00539877f
c98 110 Vss 0.00225019f
c99 109 Vss 0.00129191f
c100 101 Vss 0.00660977f
c101 92 Vss 0.00400552f
c102 83 Vss 1.70165e-19
c103 78 Vss 0.00106984f
c104 73 Vss 0.00241148f
c105 68 Vss 2.9197e-19
c106 63 Vss 0.00126608f
c107 45 Vss 0.0785271f
c108 39 Vss 0.0343198f
c109 38 Vss 0.0688517f
c110 31 Vss 7.82991e-20
c111 29 Vss 0.0338093f
c112 28 Vss 0.0998552f
c113 14 Vss 0.0835744f
c114 12 Vss 0.00226958f
c115 10 Vss 0.0837985f
c116 8 Vss 7.32238e-19
c117 6 Vss 0.0838866f
c118 4 Vss 0.0825199f
c119 2 Vss 0.00266844f
r120 141 147 0.551426
r121 141 142 13.3371
r122 140 147 0.551426
r123 139 140 4.16786
r124 135 147 0.0828784
r125 134 146 0.494161
r126 133 142 0.652036
r127 133 134 4.41793
r128 129 146 0.128424
r129 127 139 0.652036
r130 127 128 13.0037
r131 123 128 0.652036
r132 122 145 0.494161
r133 121 146 0.494161
r134 121 122 10.2946
r135 117 145 0.128424
r136 115 145 0.494161
r137 115 116 10.1279
r138 111 144 0.306046
r139 110 116 0.652036
r140 109 144 0.349767
r141 109 110 4.16786
r142 83 135 1.82344
r143 78 101 1.16709
r144 78 129 2.16729
r145 73 123 4.83471
r146 68 92 1.16709
r147 68 117 2.16729
r148 63 111 1.82344
r149 45 101 0.238214
r150 43 45 1.8672
r151 40 43 0.0685365
r152 38 43 0.5835
r153 38 39 2.8008
r154 35 39 0.652036
r155 31 92 0.238214
r156 29 31 1.45875
r157 28 32 0.652036
r158 28 31 1.45875
r159 25 29 0.652036
r160 14 40 2.5674
r161 12 83 1.16709
r162 10 35 2.5674
r163 8 73 1.16709
r164 6 32 2.5674
r165 4 25 2.5674
r166 2 63 1.16709
.ends

.subckt PM_G3_MUXI2_N1_VDD 2 4 6 8 12 14 28 38 60 62 63 66 68 72 74 75 76 77 78
+ 79 81 82 87 88 90 99 Vss
c99 99 Vss 0.00651319f
c100 90 Vss 0.00555165f
c101 88 Vss 3.54369e-19
c102 82 Vss 4.42156e-19
c103 81 Vss 0.00190072f
c104 79 Vss 0.00690705f
c105 78 Vss 8.63529e-19
c106 77 Vss 4.40622e-19
c107 76 Vss 0.00130949f
c108 75 Vss 6.09322e-19
c109 74 Vss 0.00547771f
c110 72 Vss 9.38425e-19
c111 68 Vss 0.00834424f
c112 66 Vss 0.00132511f
c113 63 Vss 6.1175e-19
c114 62 Vss 0.00344974f
c115 60 Vss 0.00121763f
c116 39 Vss 0.0805612f
c117 38 Vss 0.102888f
c118 29 Vss 0.0355046f
c119 28 Vss 0.1003f
c120 14 Vss 0.00271849f
c121 12 Vss 0.0806222f
c122 8 Vss 0.0814405f
c123 6 Vss 0.00155055f
c124 4 Vss 0.0842982f
c125 2 Vss 0.0825186f
r126 80 88 0.537385
r127 80 81 4.16786
r128 79 88 0.537385
r129 78 87 0.326018
r130 78 79 13.3788
r131 77 84 0.510562
r132 76 88 0.0936215
r133 76 77 1.35523
r134 74 87 0.326018
r135 74 75 10.1279
r136 72 99 1.16709
r137 70 75 0.652036
r138 70 72 2.16729
r139 69 82 0.494161
r140 68 81 0.652036
r141 68 69 13.0037
r142 64 82 0.128424
r143 64 66 4.83471
r144 62 82 0.494161
r145 62 63 7.46046
r146 60 90 1.16709
r147 58 63 0.652036
r148 58 60 2.16729
r149 44 99 0.238214
r150 44 46 1.92555
r151 39 46 0.5835
r152 38 40 0.652036
r153 38 39 2.8008
r154 35 46 0.0685365
r155 31 90 0.238214
r156 29 31 1.45875
r157 28 32 0.652036
r158 28 31 1.45875
r159 25 29 0.652036
r160 14 84 1.16709
r161 12 40 2.5674
r162 8 35 2.5674
r163 6 66 1.16709
r164 4 25 2.5674
r165 2 32 2.5674
.ends

.subckt PM_G3_MUXI2_N1_SELI 2 6 8 21 33 35 38 43 53 58 72 77 78 Vss
c67 78 Vss 3.71671e-19
c68 72 Vss 0.00114167f
c69 58 Vss 0.00216403f
c70 53 Vss 0.00206075f
c71 43 Vss 9.19217e-19
c72 38 Vss 0.00147194f
c73 36 Vss 0.00160147f
c74 35 Vss 0.00416276f
c75 33 Vss 0.00272744f
c76 21 Vss 0.0575023f
c77 6 Vss 0.0575023f
c78 2 Vss 0.00148239f
r79 77 78 0.655813
r80 76 77 3.501
r81 72 76 0.655813
r82 43 53 1.16709
r83 43 72 2.00578
r84 43 46 0.833571
r85 38 58 1.16709
r86 38 78 2.00578
r87 35 46 0.0685365
r88 35 36 7.46046
r89 31 36 0.652036
r90 31 33 5.58493
r91 21 58 0.50025
r92 18 53 0.50025
r93 8 21 1.80885
r94 6 18 1.80885
r95 2 33 1.16709
.ends

.subckt PM_G3_MUXI2_N1_SEL 2 4 6 8 16 22 26 36 37 40 42 46 51 58 63 68 72 77 78
+ Vss
c73 78 Vss 8.48303e-20
c74 77 Vss 2.4421e-20
c75 72 Vss 7.30413e-19
c76 68 Vss 0.00150427f
c77 63 Vss 0.00289461f
c78 58 Vss 0.00236419f
c79 51 Vss 4.10742e-19
c80 46 Vss 1.61132e-19
c81 42 Vss 0.00131501f
c82 37 Vss 0.00193143f
c83 36 Vss 6.68718e-20
c84 26 Vss 0.057622f
c85 22 Vss 0.0712295f
c86 20 Vss 0.0247918f
c87 17 Vss 0.0369263f
c88 16 Vss 0.187844f
c89 8 Vss 0.0575023f
c90 2 Vss 0.084915f
r91 76 78 0.655813
r92 76 77 3.501
r93 72 77 0.655813
r94 54 63 1.16709
r95 54 72 2.00578
r96 51 54 0.5835
r97 49 58 1.16709
r98 46 49 0.5835
r99 42 68 1.16709
r100 42 78 2.00578
r101 38 46 0.0685365
r102 38 40 1.70882
r103 37 51 0.0685365
r104 37 40 2.87582
r105 36 58 0.0476429
r106 33 68 0.50025
r107 26 63 0.50025
r108 22 58 0.357321
r109 20 36 0.326018
r110 20 22 0.40845
r111 17 36 6.7686
r112 16 36 0.326018
r113 16 36 0.1167
r114 13 17 0.652036
r115 8 33 1.80885
r116 6 26 1.80885
r117 4 22 2.15895
r118 2 13 2.5674
.ends

.subckt PM_G3_MUXI2_N1_B 2 4 7 16 20 24 27 Vss
c22 27 Vss 0.00591505f
c23 24 Vss 5.28389e-19
c24 20 Vss 0.0298499f
c25 16 Vss 0.0664813f
c26 7 Vss 0.142354f
c27 4 Vss 0.272228f
c28 2 Vss 0.0800936f
r29 24 27 1.16709
r30 16 27 0.50025
r31 16 18 1.9839
r32 12 20 0.494161
r33 9 20 0.494161
r34 8 18 0.0685365
r35 7 20 0.128424
r36 7 8 4.7847
r37 4 12 9.04425
r38 2 9 2.62575
.ends

.subckt PM_G3_MUXI2_N1_Z 2 4 30 33 Vss
c33 30 Vss 0.00283949f
c34 4 Vss 0.00148239f
c35 2 Vss 0.00156677f
r36 33 35 5.16814
r37 30 33 4.00114
r38 4 35 1.16709
r39 2 30 1.16709
.ends

.subckt PM_G3_MUXI2_N1_A 2 4 14 19 22 Vss
c24 22 Vss 0.00548526f
c25 19 Vss 4.55558e-19
c26 14 Vss 0.0830192f
c27 2 Vss 0.4453f
r28 19 22 1.16709
r29 12 22 0.238214
r30 12 14 1.92555
r31 7 14 0.0685365
r32 2 4 12.837
r33 2 7 2.5674
.ends

.subckt G3_MUXI2_N1  VSS VDD SEL B Z A
*
* A	A
* Z	Z
* B	B
* SEL	SEL
* VDD	VDD
* VSS	VSS
XI1.X0 N_SELI_XI1.X0_D N_VDD_XI1.X0_PGD N_SEL_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
XI2.X0 N_SELI_XI1.X0_D N_VSS_XI2.X0_PGD N_SEL_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_SELI_XI5.X0_CG N_B_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW1
XI3.X0 N_Z_XI3.X0_D N_VSS_XI3.X0_PGD N_SEL_XI3.X0_CG N_B_XI3.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW1
XI4.X0 N_Z_XI5.X0_D N_VDD_XI4.X0_PGD N_SEL_XI4.X0_CG N_A_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW1
XI0.X0 N_Z_XI3.X0_D N_VSS_XI0.X0_PGD N_SELI_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW1
*
x_PM_G3_MUXI2_N1_VSS N_VSS_XI1.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI5.X0_S N_VSS_XI3.X0_PGD N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_4_p
+ N_VSS_c_62_p N_VSS_c_21_p N_VSS_c_47_p N_VSS_c_5_p N_VSS_c_27_p N_VSS_c_18_p
+ N_VSS_c_29_p N_VSS_c_6_p N_VSS_c_20_p N_VSS_c_7_p N_VSS_c_11_p N_VSS_c_12_p
+ N_VSS_c_30_p N_VSS_c_25_p N_VSS_c_32_p N_VSS_c_37_p N_VSS_c_38_p VSS
+ N_VSS_c_13_p N_VSS_c_26_p N_VSS_c_39_p Vss PM_G3_MUXI2_N1_VSS
x_PM_G3_MUXI2_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI2.X0_S
+ N_VDD_XI5.X0_PGD N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_90_n N_VDD_c_181_p
+ N_VDD_c_91_n N_VDD_c_94_n N_VDD_c_100_n N_VDD_c_101_n N_VDD_c_107_n
+ N_VDD_c_113_n N_VDD_c_114_n N_VDD_c_117_n N_VDD_c_118_n N_VDD_c_119_n
+ N_VDD_c_120_n N_VDD_c_121_n N_VDD_c_126_n N_VDD_c_128_n VDD N_VDD_c_129_n
+ N_VDD_c_130_n N_VDD_c_135_p Vss PM_G3_MUXI2_N1_VDD
x_PM_G3_MUXI2_N1_SELI N_SELI_XI1.X0_D N_SELI_XI5.X0_CG N_SELI_XI0.X0_CG
+ N_SELI_c_188_n N_SELI_c_189_n N_SELI_c_192_n N_SELI_c_193_n N_SELI_c_209_n
+ N_SELI_c_211_n N_SELI_c_196_n N_SELI_c_198_n N_SELI_c_199_n N_SELI_c_231_p Vss
+ PM_G3_MUXI2_N1_SELI
x_PM_G3_MUXI2_N1_SEL N_SEL_XI1.X0_CG N_SEL_XI2.X0_CG N_SEL_XI3.X0_CG
+ N_SEL_XI4.X0_CG N_SEL_c_253_n N_SEL_c_254_n N_SEL_c_305_p N_SEL_c_255_n
+ N_SEL_c_257_n SEL N_SEL_c_258_n N_SEL_c_259_n N_SEL_c_274_n N_SEL_c_260_n
+ N_SEL_c_275_n N_SEL_c_262_n N_SEL_c_263_n N_SEL_c_265_n N_SEL_c_266_n Vss
+ PM_G3_MUXI2_N1_SEL
x_PM_G3_MUXI2_N1_B N_B_XI5.X0_PGS N_B_XI3.X0_PGS N_B_c_326_n N_B_c_344_n
+ N_B_c_336_n B N_B_c_328_n Vss PM_G3_MUXI2_N1_B
x_PM_G3_MUXI2_N1_Z N_Z_XI5.X0_D N_Z_XI3.X0_D N_Z_c_352_n Z Vss PM_G3_MUXI2_N1_Z
x_PM_G3_MUXI2_N1_A N_A_XI4.X0_PGS N_A_XI0.X0_PGS N_A_c_383_n A N_A_c_389_n Vss
+ PM_G3_MUXI2_N1_A
cc_1 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.0017188f
cc_2 N_VSS_XI3.X0_PGD N_VDD_XI5.X0_PGD 2.27468e-19
cc_3 N_VSS_XI0.X0_PGD N_VDD_XI4.X0_PGD 2.27468e-19
cc_4 N_VSS_c_4_p N_VDD_c_90_n 0.0017188f
cc_5 N_VSS_c_5_p N_VDD_c_91_n 9.32947e-19
cc_6 N_VSS_c_6_p N_VDD_c_91_n 3.82294e-19
cc_7 N_VSS_c_7_p N_VDD_c_91_n 4.10707e-19
cc_8 N_VSS_c_4_p N_VDD_c_94_n 2.72324e-19
cc_9 N_VSS_c_5_p N_VDD_c_94_n 0.00141228f
cc_10 N_VSS_c_6_p N_VDD_c_94_n 0.00112249f
cc_11 N_VSS_c_11_p N_VDD_c_94_n 0.00419135f
cc_12 N_VSS_c_12_p N_VDD_c_94_n 0.00124457f
cc_13 N_VSS_c_13_p N_VDD_c_94_n 7.74609e-19
cc_14 N_VSS_c_11_p N_VDD_c_100_n 0.00157719f
cc_15 N_VSS_XI2.X0_PGS N_VDD_c_101_n 2.93604e-19
cc_16 N_VSS_XI3.X0_PGD N_VDD_c_101_n 2.36238e-19
cc_17 N_VSS_c_5_p N_VDD_c_101_n 0.00181129f
cc_18 N_VSS_c_18_p N_VDD_c_101_n 7.45025e-19
cc_19 N_VSS_c_6_p N_VDD_c_101_n 9.55109e-19
cc_20 N_VSS_c_20_p N_VDD_c_101_n 2.60394e-19
cc_21 N_VSS_c_21_p N_VDD_c_107_n 0.00102426f
cc_22 N_VSS_c_18_p N_VDD_c_107_n 0.00161703f
cc_23 N_VSS_c_20_p N_VDD_c_107_n 2.03837e-19
cc_24 N_VSS_c_12_p N_VDD_c_107_n 0.0056811f
cc_25 N_VSS_c_25_p N_VDD_c_107_n 0.00454933f
cc_26 N_VSS_c_26_p N_VDD_c_107_n 7.61747e-19
cc_27 N_VSS_c_27_p N_VDD_c_113_n 0.00125492f
cc_28 N_VSS_XI4.X0_S N_VDD_c_114_n 3.7884e-19
cc_29 N_VSS_c_29_p N_VDD_c_114_n 4.73473e-19
cc_30 N_VSS_c_30_p N_VDD_c_114_n 0.00742779f
cc_31 N_VSS_c_30_p N_VDD_c_117_n 0.00149994f
cc_32 N_VSS_c_32_p N_VDD_c_118_n 4.31398e-19
cc_33 N_VSS_c_29_p N_VDD_c_119_n 2.14355e-19
cc_34 N_VSS_c_30_p N_VDD_c_120_n 0.00106317f
cc_35 N_VSS_XI4.X0_S N_VDD_c_121_n 9.5668e-19
cc_36 N_VSS_c_29_p N_VDD_c_121_n 0.00165395f
cc_37 N_VSS_c_37_p N_VDD_c_121_n 0.00364836f
cc_38 N_VSS_c_38_p N_VDD_c_121_n 0.0050309f
cc_39 N_VSS_c_39_p N_VDD_c_121_n 8.91588e-19
cc_40 N_VSS_c_18_p N_VDD_c_126_n 4.6996e-19
cc_41 N_VSS_c_38_p N_VDD_c_126_n 0.00295094f
cc_42 N_VSS_c_12_p N_VDD_c_128_n 0.00112088f
cc_43 N_VSS_c_38_p N_VDD_c_129_n 9.75645e-19
cc_44 N_VSS_c_5_p N_VDD_c_130_n 3.48267e-19
cc_45 N_VSS_c_6_p N_VDD_c_130_n 8.0279e-19
cc_46 N_VSS_XI1.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_47 N_VSS_c_47_p N_SELI_XI1.X0_D 3.48267e-19
cc_48 N_VSS_c_20_p N_SELI_c_188_n 0.00234241f
cc_49 N_VSS_XI1.X0_S N_SELI_c_189_n 3.48267e-19
cc_50 N_VSS_c_47_p N_SELI_c_189_n 8.47286e-19
cc_51 N_VSS_c_11_p N_SELI_c_189_n 2.65284e-19
cc_52 N_VSS_c_27_p N_SELI_c_192_n 0.00140233f
cc_53 N_VSS_c_18_p N_SELI_c_193_n 0.00135778f
cc_54 N_VSS_c_20_p N_SELI_c_193_n 4.99367e-19
cc_55 N_VSS_c_38_p N_SELI_c_193_n 9.07743e-19
cc_56 N_VSS_c_18_p N_SELI_c_196_n 4.56568e-19
cc_57 N_VSS_c_20_p N_SELI_c_196_n 0.0014909f
cc_58 N_VSS_c_30_p N_SELI_c_198_n 7.53578e-19
cc_59 N_VSS_c_38_p N_SELI_c_199_n 5.03655e-19
cc_60 N_VSS_XI2.X0_PGD N_SEL_c_253_n 4.12362e-19
cc_61 N_VSS_c_6_p N_SEL_c_254_n 0.00234241f
cc_62 N_VSS_c_62_p N_SEL_c_255_n 9.36847e-19
cc_63 N_VSS_c_6_p N_SEL_c_255_n 2.03369e-19
cc_64 N_VSS_c_12_p N_SEL_c_257_n 5.44326e-19
cc_65 N_VSS_c_38_p N_SEL_c_258_n 3.80099e-19
cc_66 N_VSS_c_5_p N_SEL_c_259_n 8.36018e-19
cc_67 N_VSS_c_5_p N_SEL_c_260_n 4.56568e-19
cc_68 N_VSS_c_6_p N_SEL_c_260_n 6.1245e-19
cc_69 N_VSS_c_20_p N_SEL_c_262_n 2.00604e-19
cc_70 N_VSS_c_12_p N_SEL_c_263_n 0.00127961f
cc_71 N_VSS_c_30_p N_SEL_c_263_n 2.81471e-19
cc_72 N_VSS_c_38_p N_SEL_c_265_n 4.36463e-19
cc_73 N_VSS_c_30_p N_SEL_c_266_n 0.00119312f
cc_74 N_VSS_XI2.X0_PGS N_B_c_326_n 2.96367e-19
cc_75 N_VSS_c_27_p B 0.00220388f
cc_76 N_VSS_XI5.X0_S N_B_c_328_n 0.00246958f
cc_77 N_VSS_c_27_p N_B_c_328_n 8.835e-19
cc_78 N_VSS_XI5.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_79 N_VSS_XI4.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_80 N_VSS_c_27_p N_Z_XI5.X0_D 3.48267e-19
cc_81 N_VSS_c_29_p N_Z_XI5.X0_D 3.48267e-19
cc_82 N_VSS_XI5.X0_S N_Z_c_352_n 3.48267e-19
cc_83 N_VSS_XI4.X0_S N_Z_c_352_n 3.48267e-19
cc_84 N_VSS_c_27_p N_Z_c_352_n 5.68449e-19
cc_85 N_VSS_c_29_p N_Z_c_352_n 5.69026e-19
cc_86 N_VSS_c_38_p N_Z_c_352_n 3.26224e-19
cc_87 N_VDD_XI2.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_88 N_VDD_c_94_n N_SELI_XI1.X0_D 3.7884e-19
cc_89 N_VDD_c_101_n N_SELI_XI1.X0_D 3.48267e-19
cc_90 N_VDD_c_135_p N_SELI_XI5.X0_CG 0.00237871f
cc_91 N_VDD_XI2.X0_S N_SELI_c_189_n 3.48267e-19
cc_92 N_VDD_c_94_n N_SELI_c_189_n 5.34437e-19
cc_93 N_VDD_c_101_n N_SELI_c_189_n 7.03427e-19
cc_94 N_VDD_c_94_n N_SELI_c_192_n 2.96638e-19
cc_95 N_VDD_c_121_n N_SELI_c_193_n 6.15494e-19
cc_96 N_VDD_c_113_n N_SELI_c_209_n 7.54639e-19
cc_97 N_VDD_c_135_p N_SELI_c_209_n 5.0614e-19
cc_98 N_VDD_c_113_n N_SELI_c_211_n 4.85469e-19
cc_99 N_VDD_c_135_p N_SELI_c_211_n 0.013665f
cc_100 N_VDD_c_121_n N_SELI_c_196_n 3.66936e-19
cc_101 N_VDD_c_130_n N_SEL_XI1.X0_CG 8.03148e-19
cc_102 N_VDD_XI1.X0_PGD N_SEL_c_253_n 4.25379e-19
cc_103 N_VDD_XI2.X0_S N_SEL_c_257_n 9.18655e-19
cc_104 N_VDD_c_101_n N_SEL_c_257_n 0.00161606f
cc_105 N_VDD_c_107_n N_SEL_c_258_n 2.90143e-19
cc_106 N_VDD_c_114_n N_SEL_c_258_n 3.06021e-19
cc_107 N_VDD_c_121_n N_SEL_c_258_n 6.68274e-19
cc_108 N_VDD_c_107_n N_SEL_c_274_n 2.1079e-19
cc_109 N_VDD_c_107_n N_SEL_c_275_n 2.19082e-19
cc_110 N_VDD_c_135_p N_SEL_c_275_n 2.00604e-19
cc_111 N_VDD_XI4.X0_PGD N_SEL_c_262_n 3.11814e-19
cc_112 N_VDD_c_121_n N_SEL_c_262_n 3.66936e-19
cc_113 N_VDD_c_107_n N_SEL_c_263_n 4.86613e-19
cc_114 N_VDD_c_121_n N_SEL_c_265_n 2.2501e-19
cc_115 N_VDD_c_114_n N_Z_XI5.X0_D 3.7884e-19
cc_116 N_VDD_XI2.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_117 N_VDD_XI0.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_118 N_VDD_c_101_n N_Z_XI3.X0_D 3.48267e-19
cc_119 N_VDD_c_107_n N_Z_XI3.X0_D 3.7884e-19
cc_120 N_VDD_c_119_n N_Z_XI3.X0_D 3.72199e-19
cc_121 N_VDD_XI2.X0_S N_Z_c_352_n 3.48267e-19
cc_122 N_VDD_XI0.X0_S N_Z_c_352_n 3.48267e-19
cc_123 N_VDD_c_101_n N_Z_c_352_n 8.10024e-19
cc_124 N_VDD_c_107_n N_Z_c_352_n 5.35804e-19
cc_125 N_VDD_c_114_n N_Z_c_352_n 5.35804e-19
cc_126 N_VDD_c_119_n N_Z_c_352_n 8.05266e-19
cc_127 N_VDD_c_121_n N_Z_c_352_n 7.45211e-19
cc_128 N_VDD_XI4.X0_PGD N_A_XI4.X0_PGS 0.00162178f
cc_129 N_VDD_c_121_n N_A_XI4.X0_PGS 0.0010699f
cc_130 N_VDD_c_114_n N_A_c_383_n 3.3974e-19
cc_131 N_VDD_c_121_n N_A_c_383_n 4.15738e-19
cc_132 N_VDD_c_113_n A 5.43314e-19
cc_133 N_VDD_c_114_n A 0.00141439f
cc_134 N_VDD_c_121_n A 5.04211e-19
cc_135 N_VDD_c_135_p A 3.48267e-19
cc_136 N_VDD_c_181_p N_A_c_389_n 0.00480616f
cc_137 N_VDD_c_113_n N_A_c_389_n 3.89161e-19
cc_138 N_VDD_c_114_n N_A_c_389_n 0.00117371f
cc_139 N_VDD_c_121_n N_A_c_389_n 4.41003e-19
cc_140 N_VDD_c_135_p N_A_c_389_n 6.39485e-19
cc_141 N_SELI_c_189_n N_SEL_c_253_n 8.93041e-19
cc_142 N_SELI_c_192_n N_SEL_c_253_n 3.46631e-19
cc_143 N_SELI_c_209_n N_SEL_c_257_n 0.00339809f
cc_144 N_SELI_c_193_n N_SEL_c_258_n 0.00240446f
cc_145 N_SELI_c_189_n N_SEL_c_259_n 0.0021504f
cc_146 N_SELI_c_192_n N_SEL_c_259_n 0.00339809f
cc_147 N_SELI_c_189_n N_SEL_c_260_n 9.71051e-19
cc_148 N_SELI_c_192_n N_SEL_c_260_n 6.41327e-19
cc_149 N_SELI_c_209_n N_SEL_c_275_n 7.09664e-19
cc_150 N_SELI_c_211_n N_SEL_c_275_n 0.00496695f
cc_151 N_SELI_c_196_n N_SEL_c_275_n 8.74049e-19
cc_152 N_SELI_c_193_n N_SEL_c_262_n 4.99367e-19
cc_153 N_SELI_c_211_n N_SEL_c_262_n 8.86313e-19
cc_154 N_SELI_c_196_n N_SEL_c_262_n 0.00491002f
cc_155 N_SELI_c_193_n N_SEL_c_263_n 0.00165721f
cc_156 N_SELI_c_209_n N_SEL_c_263_n 4.70859e-19
cc_157 N_SELI_c_198_n N_SEL_c_263_n 9.36901e-19
cc_158 N_SELI_c_231_p N_SEL_c_263_n 7.85443e-19
cc_159 N_SELI_c_189_n N_SEL_c_265_n 2.46723e-19
cc_160 N_SELI_c_209_n N_SEL_c_265_n 2.46502e-19
cc_161 N_SELI_c_199_n N_SEL_c_265_n 0.00142585f
cc_162 N_SELI_c_209_n N_SEL_c_266_n 0.00166116f
cc_163 N_SELI_c_198_n N_SEL_c_266_n 7.57935e-19
cc_164 N_SELI_XI5.X0_CG N_B_XI5.X0_PGS 4.34645e-19
cc_165 N_SELI_c_211_n N_B_XI5.X0_PGS 6.90642e-19
cc_166 N_SELI_c_189_n N_B_XI3.X0_PGS 2.37944e-19
cc_167 N_SELI_c_192_n N_B_XI3.X0_PGS 3.60699e-19
cc_168 N_SELI_c_211_n N_B_XI3.X0_PGS 5.45575e-19
cc_169 N_SELI_c_192_n N_B_c_326_n 3.87281e-19
cc_170 N_SELI_c_192_n N_B_c_336_n 5.40503e-19
cc_171 N_SELI_c_192_n B 0.0012892f
cc_172 N_SELI_c_192_n N_B_c_328_n 0.00106294f
cc_173 N_SELI_c_189_n N_Z_c_352_n 5.41397e-19
cc_174 N_SELI_c_193_n N_Z_c_352_n 0.00205681f
cc_175 N_SELI_c_209_n N_Z_c_352_n 0.00246976f
cc_176 N_SELI_c_211_n N_Z_c_352_n 9.16045e-19
cc_177 N_SELI_c_188_n N_A_XI4.X0_PGS 4.5346e-19
cc_178 N_SELI_c_196_n N_A_XI4.X0_PGS 0.00276355f
cc_179 N_SELI_c_196_n N_A_c_389_n 2.00604e-19
cc_180 N_SEL_c_254_n N_B_XI3.X0_PGS 2.04953e-19
cc_181 N_SEL_c_305_p N_B_XI3.X0_PGS 4.64062e-19
cc_182 N_SEL_c_257_n N_B_XI3.X0_PGS 8.04174e-19
cc_183 N_SEL_c_260_n N_B_XI3.X0_PGS 0.00100354f
cc_184 N_SEL_c_275_n N_B_XI3.X0_PGS 0.00142122f
cc_185 N_SEL_c_257_n N_B_c_344_n 2.97958e-19
cc_186 N_SEL_c_260_n N_B_c_344_n 3.50453e-19
cc_187 N_SEL_c_260_n N_B_c_328_n 9.99041e-19
cc_188 N_SEL_c_258_n N_Z_c_352_n 0.00187327f
cc_189 N_SEL_c_274_n N_Z_c_352_n 0.00194252f
cc_190 N_SEL_c_275_n N_Z_c_352_n 9.12105e-19
cc_191 N_SEL_c_262_n N_Z_c_352_n 9.02042e-19
cc_192 N_SEL_c_263_n N_Z_c_352_n 8.60225e-19
cc_193 N_SEL_c_265_n N_Z_c_352_n 0.0021646f
cc_194 N_SEL_c_266_n N_Z_c_352_n 8.38981e-19
cc_195 N_SEL_XI4.X0_CG N_A_XI4.X0_PGS 4.42555e-19
cc_196 N_SEL_c_262_n N_A_XI4.X0_PGS 0.00276355f
cc_197 N_SEL_c_258_n A 7.0885e-19
cc_198 N_SEL_c_262_n A 4.56568e-19
cc_199 N_SEL_XI4.X0_CG N_A_c_389_n 0.00234241f
cc_200 N_SEL_c_258_n N_A_c_389_n 4.99367e-19
cc_201 N_SEL_c_262_n N_A_c_389_n 0.0014909f
cc_202 N_B_XI5.X0_PGS N_A_XI4.X0_PGS 0.00137535f
*
.ends
*
*
.subckt MUXI2_HPNW1 A B S0 Y VDD VSS
xgate (VSS VDD S0 B Y A) G3_MUXI2_N1
.ends
*
* File: G2_NAND2_N1.pex.netlist
* Created: Tue Feb 22 16:31:07 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NAND2_N1_VSS 2 4 6 8 10 20 23 45 50 59 68 69 70 Vss
c27 70 Vss 7.84263e-19
c28 69 Vss 0.00114439f
c29 59 Vss 0.00441797f
c30 50 Vss 5.92201e-19
c31 45 Vss 0.00559837f
c32 38 Vss 0.0299355f
c33 37 Vss 0.0299355f
c34 32 Vss 0.105919f
c35 27 Vss 0.0688517f
c36 23 Vss 6.52493e-20
c37 21 Vss 0.0348456f
c38 20 Vss 0.064644f
c39 10 Vss 0.0834601f
c40 8 Vss 0.0831275f
c41 6 Vss 0.0830428f
c42 4 Vss 0.0828837f
c43 2 Vss 0.00278021f
r44 69 71 0.652036
r45 69 70 1.66714
r46 63 70 0.652036
r47 63 68 9.12761
r48 50 59 1.16709
r49 50 71 2.16729
r50 45 68 4.87639
r51 33 38 0.494161
r52 32 34 0.652036
r53 32 33 2.9175
r54 29 38 0.128424
r55 28 37 0.494161
r56 27 38 0.494161
r57 27 28 2.8008
r58 24 37 0.128424
r59 23 59 0.238214
r60 21 23 1.4004
r61 20 37 0.494161
r62 20 23 1.5171
r63 17 21 0.652036
r64 10 34 2.5674
r65 8 29 2.5674
r66 6 17 2.5674
r67 4 24 2.5674
r68 2 45 1.16709
.ends

.subckt PM_G2_NAND2_N1_VDD 2 4 6 15 17 31 33 34 35 42 44 50 Vss
c43 50 Vss 0.00511687f
c44 42 Vss 0.00686567f
c45 40 Vss 0.00174586f
c46 35 Vss 0.00426091f
c47 34 Vss 8.36616e-19
c48 33 Vss 0.00735566f
c49 31 Vss 0.00189708f
c50 17 Vss 0.184529f
c51 15 Vss 0.0364084f
c52 6 Vss 0.00252742f
c53 4 Vss 0.00226556f
c54 2 Vss 0.0989662f
r55 40 44 0.326018
r56 40 42 4.83471
r57 39 42 7.002
r58 37 50 1.16709
r59 35 39 0.655813
r60 35 37 2.04225
r61 33 44 0.326018
r62 33 34 10.3363
r63 29 34 0.652036
r64 29 31 4.83471
r65 17 50 0.50025
r66 15 17 5.11257
r67 12 15 0.652541
r68 6 42 1.16709
r69 4 31 1.16709
r70 2 12 3.2676
.ends

.subckt PM_G2_NAND2_N1_A 2 4 13 18 21 26 31 Vss
c21 31 Vss 0.00366686f
c22 26 Vss 0.00318863f
c23 18 Vss 0.00132825f
c24 13 Vss 0.0578401f
c25 2 Vss 0.0573541f
r26 23 31 1.16709
r27 21 23 1.91721
r28 18 26 1.16709
r29 18 21 2.9175
r30 13 31 0.50025
r31 10 26 0.50025
r32 4 13 1.80885
r33 2 10 1.80885
.ends

.subckt PM_G2_NAND2_N1_Z 2 4 25 28 Vss
c25 25 Vss 0.00107312f
c26 4 Vss 0.00148239f
c27 2 Vss 0.00149062f
r28 28 30 4.58464
r29 25 28 4.58464
r30 4 30 1.16709
r31 2 25 1.16709
.ends

.subckt PM_G2_NAND2_N1_B 2 4 10 11 14 18 21 Vss
c24 18 Vss 1.08854e-19
c25 14 Vss 0.147604f
c26 11 Vss 0.0356774f
c27 10 Vss 0.286243f
c28 2 Vss 0.174968f
r29 18 21 0.0416786
r30 14 18 1.16709
r31 12 14 2.8008
r32 10 12 0.652036
r33 10 11 8.92755
r34 7 11 0.652036
r35 4 14 3.0342
r36 2 7 5.835
.ends

.subckt G2_NAND2_N1  VSS VDD A Z B
*
* B	B
* Z	Z
* A	A
* VDD	VDD
* VSS	VSS
XI7.X0 N_Z_XI7.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_B_XI7.X0_PGS N_VSS_XI7.X0_S
+ TIGFET_HPNW1
XI8.X0 N_Z_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW1
XI9.X0 N_Z_XI8.X0_D N_VSS_XI9.X0_PGD N_B_XI9.X0_CG N_VSS_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW1
*
x_PM_G2_NAND2_N1_VSS N_VSS_XI7.X0_S N_VSS_XI8.X0_PGD N_VSS_XI8.X0_PGS
+ N_VSS_XI9.X0_PGD N_VSS_XI9.X0_PGS N_VSS_c_6_p N_VSS_c_18_p N_VSS_c_1_p
+ N_VSS_c_4_p N_VSS_c_5_p VSS N_VSS_c_9_p N_VSS_c_10_p Vss PM_G2_NAND2_N1_VSS
x_PM_G2_NAND2_N1_VDD N_VDD_XI7.X0_PGD N_VDD_XI8.X0_S N_VDD_XI9.X0_S N_VDD_c_61_p
+ N_VDD_c_54_p N_VDD_c_29_n N_VDD_c_33_n N_VDD_c_37_n N_VDD_c_57_p N_VDD_c_38_n
+ VDD N_VDD_c_43_p Vss PM_G2_NAND2_N1_VDD
x_PM_G2_NAND2_N1_A N_A_XI7.X0_CG N_A_XI8.X0_CG N_A_c_71_n N_A_c_72_n A
+ N_A_c_79_n N_A_c_75_n Vss PM_G2_NAND2_N1_A
x_PM_G2_NAND2_N1_Z N_Z_XI7.X0_D N_Z_XI8.X0_D N_Z_c_94_n Z Vss PM_G2_NAND2_N1_Z
x_PM_G2_NAND2_N1_B N_B_XI7.X0_PGS N_B_XI9.X0_CG N_B_c_117_n N_B_c_119_n
+ N_B_c_123_n N_B_c_127_n B Vss PM_G2_NAND2_N1_B
cc_1 N_VSS_c_1_p N_VDD_XI8.X0_S 0.00136022f
cc_2 N_VSS_XI8.X0_PGS N_VDD_c_29_n 4.05134e-19
cc_3 N_VSS_c_1_p N_VDD_c_29_n 0.00385472f
cc_4 N_VSS_c_4_p N_VDD_c_29_n 0.00232594f
cc_5 N_VSS_c_5_p N_VDD_c_29_n 0.00101015f
cc_6 N_VSS_c_6_p N_VDD_c_33_n 0.00171596f
cc_7 N_VSS_c_4_p N_VDD_c_33_n 0.00161703f
cc_8 N_VSS_c_5_p N_VDD_c_33_n 2.03837e-19
cc_9 N_VSS_c_9_p N_VDD_c_33_n 0.00286543f
cc_10 N_VSS_c_10_p N_VDD_c_37_n 0.00103397f
cc_11 N_VSS_XI9.X0_PGS N_VDD_c_38_n 4.47716e-19
cc_12 N_VSS_c_1_p N_VDD_c_38_n 2.23518e-19
cc_13 N_VSS_c_4_p N_VDD_c_38_n 5.24284e-19
cc_14 N_VSS_c_5_p N_A_c_71_n 0.00234241f
cc_15 N_VSS_c_1_p N_A_c_72_n 0.00297841f
cc_16 N_VSS_c_4_p N_A_c_72_n 8.12473e-19
cc_17 N_VSS_c_5_p N_A_c_72_n 5.42695e-19
cc_18 N_VSS_c_18_p N_A_c_75_n 7.84334e-19
cc_19 N_VSS_c_4_p N_A_c_75_n 4.56568e-19
cc_20 N_VSS_c_5_p N_A_c_75_n 0.00184767f
cc_21 N_VSS_XI7.X0_S N_Z_XI7.X0_D 3.43419e-19
cc_22 N_VSS_c_1_p N_Z_XI7.X0_D 3.48267e-19
cc_23 N_VSS_XI7.X0_S N_Z_c_94_n 3.48267e-19
cc_24 N_VSS_c_1_p N_Z_c_94_n 0.00178967f
cc_25 N_VSS_XI8.X0_PGD N_B_c_117_n 6.72196e-19
cc_26 N_VSS_XI9.X0_PGD N_B_c_117_n 6.72196e-19
cc_27 N_VSS_XI8.X0_PGS N_B_c_119_n 7.91098e-19
cc_28 N_VDD_XI7.X0_PGD N_A_XI7.X0_CG 4.91184e-19
cc_29 N_VDD_XI7.X0_PGD N_A_c_79_n 2.88617e-19
cc_30 N_VDD_c_43_p N_A_c_79_n 7.96439e-19
cc_31 N_VDD_c_33_n N_A_c_75_n 2.29043e-19
cc_32 N_VDD_c_43_p N_Z_XI7.X0_D 0.00132057f
cc_33 N_VDD_XI8.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_34 N_VDD_XI9.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_35 N_VDD_c_29_n N_Z_XI8.X0_D 3.48267e-19
cc_36 N_VDD_c_33_n N_Z_XI8.X0_D 3.7884e-19
cc_37 N_VDD_c_38_n N_Z_XI8.X0_D 3.48267e-19
cc_38 N_VDD_XI7.X0_PGD N_Z_c_94_n 3.00781e-19
cc_39 N_VDD_XI8.X0_S N_Z_c_94_n 3.48267e-19
cc_40 N_VDD_XI9.X0_S N_Z_c_94_n 3.48267e-19
cc_41 N_VDD_c_54_p N_Z_c_94_n 7.07078e-19
cc_42 N_VDD_c_29_n N_Z_c_94_n 5.69026e-19
cc_43 N_VDD_c_33_n N_Z_c_94_n 7.07375e-19
cc_44 N_VDD_c_57_p N_Z_c_94_n 0.00174191f
cc_45 N_VDD_c_38_n N_Z_c_94_n 0.00291831f
cc_46 N_VDD_c_43_p N_Z_c_94_n 8.835e-19
cc_47 N_VDD_XI7.X0_PGD N_B_XI7.X0_PGS 0.00320747f
cc_48 N_VDD_c_61_p N_B_c_117_n 0.0097987f
cc_49 N_VDD_c_38_n N_B_c_117_n 2.48119e-19
cc_50 N_VDD_c_33_n N_B_c_123_n 4.73957e-19
cc_51 N_VDD_c_57_p N_B_c_123_n 3.81676e-19
cc_52 N_VDD_c_38_n N_B_c_123_n 0.001001f
cc_53 N_VDD_c_43_p N_B_c_123_n 0.00150149f
cc_54 N_VDD_c_33_n N_B_c_127_n 4.10393e-19
cc_55 N_VDD_c_57_p N_B_c_127_n 5.19718e-19
cc_56 N_VDD_c_38_n N_B_c_127_n 0.00144738f
cc_57 N_VDD_c_43_p N_B_c_127_n 3.81676e-19
cc_58 N_A_c_72_n N_Z_c_94_n 0.00754545f
cc_59 N_A_c_79_n N_Z_c_94_n 9.58524e-19
cc_60 N_A_c_75_n N_Z_c_94_n 9.18163e-19
cc_61 N_A_XI7.X0_CG N_B_XI7.X0_PGS 4.5346e-19
cc_62 N_A_c_72_n N_B_XI7.X0_PGS 2.82086e-19
cc_63 N_A_c_79_n N_B_XI7.X0_PGS 5.70584e-19
cc_64 N_A_c_72_n N_B_c_117_n 3.21972e-19
cc_65 N_A_c_79_n N_B_c_117_n 0.0014179f
cc_66 N_A_c_75_n N_B_c_117_n 0.00112482f
cc_67 N_A_c_75_n N_B_c_123_n 9.27569e-19
cc_68 N_Z_c_94_n N_B_c_117_n 3.90525e-19
cc_69 N_Z_c_94_n N_B_c_123_n 9.49424e-19
cc_70 N_Z_c_94_n N_B_c_127_n 0.00147334f
*
.ends
*
*
.subckt NAND2_HPNW1 A B Y VDD VSS
xgate (VSS VDD A Y B) G2_NAND2_N1
.ends
*
* File: G2_NOR2_N1.pex.netlist
* Created: Mon Feb 28 09:28:35 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NOR2_N1_VSS 2 4 6 16 18 31 36 41 50 61 62 66 67 72 79 80 Vss
c43 80 Vss 3.75522e-19
c44 79 Vss 0.00223955f
c45 74 Vss 0.00269784f
c46 72 Vss 0.00694708f
c47 67 Vss 8.20725e-19
c48 66 Vss 0.00177669f
c49 62 Vss 6.45375e-19
c50 61 Vss 0.00385292f
c51 50 Vss 0.00491203f
c52 41 Vss 7.10513e-22
c53 36 Vss 9.27479e-19
c54 31 Vss 0.00114656f
c55 18 Vss 0.0881492f
c56 16 Vss 6.95992e-20
c57 6 Vss 0.00202759f
c58 4 Vss 0.0834348f
c59 2 Vss 0.00226843f
r60 78 79 4.16786
r61 74 78 0.655813
r62 73 80 0.494161
r63 72 79 0.652036
r64 72 73 10.1279
r65 68 80 0.128424
r66 66 80 0.494161
r67 66 67 4.37625
r68 59 67 0.652036
r69 59 61 8.46075
r70 58 62 0.655813
r71 58 61 4.87639
r72 41 74 1.82344
r73 36 50 1.16709
r74 36 68 2.16729
r75 31 62 1.82344
r76 16 50 0.238214
r77 16 18 2.04225
r78 12 18 0.0685365
r79 6 41 1.16709
r80 4 12 2.5674
r81 2 31 1.16709
.ends

.subckt PM_G2_NOR2_N1_VDD 2 4 6 8 10 27 29 45 47 48 52 54 55 57 60 64 66 72 78
+ Vss
c51 78 Vss 0.0058262f
c52 72 Vss 0.00492692f
c53 66 Vss 3.56526e-19
c54 64 Vss 9.96234e-19
c55 60 Vss 0.00134431f
c56 55 Vss 8.63545e-19
c57 54 Vss 0.0060792f
c58 52 Vss 0.0016605f
c59 49 Vss 0.00173366f
c60 48 Vss 0.00489508f
c61 47 Vss 0.00194735f
c62 45 Vss 0.00746951f
c63 37 Vss 0.127438f
c64 29 Vss 7.35265e-20
c65 27 Vss 0.0346129f
c66 26 Vss 0.101192f
c67 10 Vss 0.0842957f
c68 8 Vss 0.0823812f
c69 6 Vss 0.00220559f
c70 4 Vss 0.0830779f
c71 2 Vss 0.0842392f
r72 72 75 0.05
r73 64 78 1.16709
r74 62 64 2.16729
r75 60 75 1.16709
r76 58 60 2.20896
r77 55 57 9.04425
r78 54 62 0.652036
r79 54 57 1.12532
r80 50 66 0.0828784
r81 50 52 1.82344
r82 48 58 0.652036
r83 48 49 4.37625
r84 47 55 0.652036
r85 46 66 0.551426
r86 46 47 4.16786
r87 45 66 0.551426
r88 44 49 0.652036
r89 44 45 13.3371
r90 36 72 0.262036
r91 36 37 2.26917
r92 33 36 2.26917
r93 29 78 0.238214
r94 27 29 1.5171
r95 26 30 0.652036
r96 26 29 1.4004
r97 23 27 0.652036
r98 20 37 0.00605528
r99 17 33 0.00605528
r100 10 30 2.5674
r101 8 23 2.5674
r102 6 52 1.16709
r103 4 17 2.5674
r104 2 20 2.5674
.ends

.subckt PM_G2_NOR2_N1_B 2 4 10 13 18 21 26 31 Vss
c25 31 Vss 0.00183593f
c26 26 Vss 0.00362926f
c27 18 Vss 9.68961e-19
c28 13 Vss 0.057478f
c29 10 Vss 6.74849e-20
c30 2 Vss 0.0576626f
r31 23 31 1.16709
r32 21 23 2.20896
r33 18 26 1.16709
r34 18 21 2.62575
r35 13 31 0.50025
r36 10 26 0.50025
r37 4 13 1.80885
r38 2 10 1.80885
.ends

.subckt PM_G2_NOR2_N1_Z 2 4 25 28 Vss
c21 25 Vss 0.00301088f
c22 4 Vss 0.00148239f
c23 2 Vss 0.0021264f
r24 28 30 3.12589
r25 25 28 6.04339
r26 4 30 1.16709
r27 2 25 1.16709
.ends

.subckt PM_G2_NOR2_N1_A 2 4 10 11 14 20 Vss
c18 20 Vss 2.48297e-19
c19 14 Vss 0.116468f
c20 11 Vss 0.0348164f
c21 10 Vss 0.273262f
c22 2 Vss 0.14291f
r23 20 26 1.16709
r24 14 26 0.05
r25 12 14 1.6338
r26 10 12 0.652036
r27 10 11 8.92755
r28 7 11 0.652036
r29 4 14 3.0342
r30 2 7 4.668
.ends

.subckt G2_NOR2_N1  VSS VDD B Z A
*
* A	A
* Z	Z
* B	B
* VDD	VDD
* VSS	VSS
XI2.X0 N_Z_XI2.X0_D N_VDD_XI2.X0_PGD N_B_XI2.X0_CG N_VDD_XI2.X0_PGS
+ N_VSS_XI2.X0_S TIGFET_HPNW1
XI0.X0 N_Z_XI0.X0_D N_VSS_XI0.X0_PGD N_B_XI0.X0_CG N_A_XI0.X0_PGS N_VDD_XI0.X0_S
+ TIGFET_HPNW1
XI1.X0 N_Z_XI0.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
*
x_PM_G2_NOR2_N1_VSS N_VSS_XI2.X0_S N_VSS_XI0.X0_PGD N_VSS_XI1.X0_S N_VSS_c_31_p
+ N_VSS_c_2_p N_VSS_c_4_p N_VSS_c_7_p N_VSS_c_37_p N_VSS_c_8_p VSS N_VSS_c_6_p
+ N_VSS_c_16_p N_VSS_c_19_p N_VSS_c_17_p N_VSS_c_22_p N_VSS_c_18_p Vss
+ PM_G2_NOR2_N1_VSS
x_PM_G2_NOR2_N1_VDD N_VDD_XI2.X0_PGD N_VDD_XI2.X0_PGS N_VDD_XI0.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_c_45_n N_VDD_c_90_p N_VDD_c_46_n
+ N_VDD_c_50_n N_VDD_c_53_n N_VDD_c_55_n N_VDD_c_56_n N_VDD_c_62_n VDD
+ N_VDD_c_72_p N_VDD_c_63_n N_VDD_c_66_n N_VDD_c_69_p N_VDD_c_67_n Vss
+ PM_G2_NOR2_N1_VDD
x_PM_G2_NOR2_N1_B N_B_XI2.X0_CG N_B_XI0.X0_CG N_B_c_104_n N_B_c_95_n N_B_c_96_n
+ B N_B_c_99_n N_B_c_100_n Vss PM_G2_NOR2_N1_B
x_PM_G2_NOR2_N1_Z N_Z_XI2.X0_D N_Z_XI0.X0_D N_Z_c_124_n Z Vss PM_G2_NOR2_N1_Z
x_PM_G2_NOR2_N1_A N_A_XI0.X0_PGS N_A_XI1.X0_CG N_A_c_141_n N_A_c_145_n
+ N_A_c_147_n A Vss PM_G2_NOR2_N1_A
cc_1 N_VSS_XI0.X0_PGD N_VDD_XI1.X0_PGD 0.00180308f
cc_2 N_VSS_c_2_p N_VDD_c_45_n 0.00180308f
cc_3 N_VSS_XI2.X0_S N_VDD_c_46_n 9.5668e-19
cc_4 N_VSS_c_4_p N_VDD_c_46_n 0.00165395f
cc_5 VSS N_VDD_c_46_n 0.00476397f
cc_6 N_VSS_c_6_p N_VDD_c_46_n 0.00186257f
cc_7 N_VSS_c_7_p N_VDD_c_50_n 4.43871e-19
cc_8 N_VSS_c_8_p N_VDD_c_50_n 3.66936e-19
cc_9 VSS N_VDD_c_50_n 0.00285866f
cc_10 N_VSS_XI2.X0_S N_VDD_c_53_n 3.7884e-19
cc_11 N_VSS_c_4_p N_VDD_c_53_n 0.00104703f
cc_12 N_VSS_c_4_p N_VDD_c_55_n 7.47067e-19
cc_13 N_VSS_c_2_p N_VDD_c_56_n 3.37151e-19
cc_14 N_VSS_c_7_p N_VDD_c_56_n 0.00141228f
cc_15 N_VSS_c_8_p N_VDD_c_56_n 0.00112249f
cc_16 N_VSS_c_16_p N_VDD_c_56_n 0.0034844f
cc_17 N_VSS_c_17_p N_VDD_c_56_n 0.00588723f
cc_18 N_VSS_c_18_p N_VDD_c_56_n 7.74609e-19
cc_19 N_VSS_c_19_p N_VDD_c_62_n 0.00106075f
cc_20 N_VSS_c_7_p N_VDD_c_63_n 0.00106112f
cc_21 N_VSS_c_8_p N_VDD_c_63_n 3.95933e-19
cc_22 N_VSS_c_22_p N_VDD_c_63_n 3.86251e-19
cc_23 VSS N_VDD_c_66_n 0.00116512f
cc_24 N_VSS_c_7_p N_VDD_c_67_n 3.44698e-19
cc_25 N_VSS_c_8_p N_VDD_c_67_n 7.95135e-19
cc_26 N_VSS_c_8_p N_B_c_95_n 0.00234321f
cc_27 N_VSS_c_7_p N_B_c_96_n 8.39582e-19
cc_28 N_VSS_c_8_p N_B_c_96_n 5.42695e-19
cc_29 VSS N_B_c_96_n 0.00148607f
cc_30 N_VSS_c_8_p N_B_c_99_n 2.00604e-19
cc_31 N_VSS_c_31_p N_B_c_100_n 8.37306e-19
cc_32 N_VSS_c_7_p N_B_c_100_n 4.56568e-19
cc_33 N_VSS_c_8_p N_B_c_100_n 0.00173573f
cc_34 N_VSS_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_35 N_VSS_c_4_p N_Z_XI2.X0_D 3.48267e-19
cc_36 N_VSS_XI1.X0_S N_Z_XI0.X0_D 3.43419e-19
cc_37 N_VSS_c_37_p N_Z_XI0.X0_D 3.48267e-19
cc_38 N_VSS_c_4_p N_Z_c_124_n 8.89782e-19
cc_39 N_VSS_c_37_p N_Z_c_124_n 6.0686e-19
cc_40 VSS N_Z_c_124_n 4.63431e-19
cc_41 N_VSS_c_17_p N_Z_c_124_n 2.55365e-19
cc_42 N_VSS_XI0.X0_PGD N_A_c_141_n 9.39677e-19
cc_43 N_VSS_c_2_p N_A_c_141_n 2.16729e-19
cc_44 N_VDD_c_69_p N_B_XI2.X0_CG 0.00237871f
cc_45 N_VDD_c_69_p N_B_c_104_n 0.0010681f
cc_46 N_VDD_c_46_n N_B_c_96_n 0.0025037f
cc_47 N_VDD_c_72_p N_B_c_96_n 7.41679e-19
cc_48 N_VDD_c_69_p N_B_c_96_n 5.48133e-19
cc_49 N_VDD_c_46_n N_B_c_99_n 4.9897e-19
cc_50 N_VDD_c_72_p N_B_c_99_n 4.91501e-19
cc_51 N_VDD_c_69_p N_B_c_99_n 0.00150793f
cc_52 N_VDD_c_46_n N_B_c_100_n 3.66936e-19
cc_53 N_VDD_c_69_p N_B_c_100_n 2.00604e-19
cc_54 N_VDD_XI0.X0_S N_Z_XI0.X0_D 3.43419e-19
cc_55 N_VDD_c_55_n N_Z_XI0.X0_D 3.72199e-19
cc_56 N_VDD_c_56_n N_Z_XI0.X0_D 3.7884e-19
cc_57 N_VDD_XI0.X0_S N_Z_c_124_n 3.48267e-19
cc_58 N_VDD_c_46_n N_Z_c_124_n 5.1034e-19
cc_59 N_VDD_c_55_n N_Z_c_124_n 7.89245e-19
cc_60 N_VDD_c_56_n N_Z_c_124_n 5.36364e-19
cc_61 N_VDD_XI2.X0_PGD N_A_c_141_n 5.10213e-19
cc_62 N_VDD_XI1.X0_PGD N_A_c_141_n 2.48727e-19
cc_63 N_VDD_XI2.X0_PGS N_A_c_145_n 6.4837e-19
cc_64 N_VDD_c_46_n N_A_c_145_n 3.16598e-19
cc_65 N_VDD_c_90_p N_A_c_147_n 8.9931e-19
cc_66 N_VDD_c_63_n N_A_c_147_n 4.91217e-19
cc_67 N_VDD_c_67_n N_A_c_147_n 0.00320668f
cc_68 N_VDD_c_63_n A 6.1931e-19
cc_69 N_VDD_c_67_n A 4.56568e-19
cc_70 N_B_c_96_n N_Z_c_124_n 0.00744925f
cc_71 N_B_c_99_n N_Z_c_124_n 9.58524e-19
cc_72 N_B_c_100_n N_Z_c_124_n 8.92526e-19
cc_73 N_B_c_95_n N_A_XI0.X0_PGS 4.5346e-19
cc_74 N_B_c_100_n N_A_XI0.X0_PGS 7.86826e-19
cc_75 N_B_c_99_n N_A_c_141_n 9.25308e-19
cc_76 N_B_c_100_n N_A_c_147_n 7.50183e-19
cc_77 N_Z_c_124_n N_A_c_141_n 9.72643e-19
cc_78 N_Z_c_124_n N_A_c_147_n 9.67259e-19
cc_79 N_Z_c_124_n A 0.00155484f
*
.ends
*
*
.subckt NOR2_HPNW1 A B Y VDD VSS
xgate (VSS VDD B Y A) G2_NOR2_N1
.ends
*
* File: G2_OAI21_N1.pex.netlist
* Created: Wed Feb 23 15:42:41 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_OAI21_N1_VSS 2 4 6 8 10 22 29 45 50 55 64 73 74 78 84 86 91 94 Vss
c49 92 Vss 5.73928e-19
c50 91 Vss 0.00675279f
c51 86 Vss 0.00175471f
c52 84 Vss 0.00280649f
c53 79 Vss 0.00136179f
c54 78 Vss 0.00706512f
c55 74 Vss 6.45375e-19
c56 73 Vss 0.00483551f
c57 64 Vss 0.00536833f
c58 55 Vss 1.70165e-19
c59 50 Vss 0.00185649f
c60 45 Vss 0.0012795f
c61 33 Vss 0.0307391f
c62 29 Vss 7.39492e-20
c63 26 Vss 0.101218f
c64 22 Vss 0.0345446f
c65 21 Vss 0.0712517f
c66 10 Vss 0.0820743f
c67 8 Vss 0.0810902f
c68 6 Vss 0.00226958f
c69 4 Vss 0.0806996f
c70 2 Vss 0.00266945f
r71 91 94 0.326018
r72 90 91 13.3371
r73 86 90 0.655813
r74 85 92 0.494161
r75 84 94 0.326018
r76 84 85 4.33457
r77 80 92 0.128424
r78 78 92 0.494161
r79 78 79 10.1696
r80 73 79 0.652036
r81 72 74 0.655813
r82 72 73 13.3371
r83 55 86 1.82344
r84 50 64 1.16709
r85 50 80 2.16729
r86 45 74 1.82344
r87 29 64 0.238214
r88 27 33 0.494161
r89 27 29 1.5171
r90 26 30 0.652036
r91 26 29 1.4004
r92 23 33 0.128424
r93 21 33 0.494161
r94 21 22 2.8008
r95 18 22 0.652036
r96 10 30 2.5674
r97 8 23 2.5674
r98 6 55 1.16709
r99 4 18 2.5674
r100 2 45 1.16709
.ends

.subckt PM_G2_OAI21_N1_VDD 2 4 6 8 38 39 41 43 47 49 51 56 59 65 Vss
c51 65 Vss 0.00591189f
c52 57 Vss 5.34798e-19
c53 56 Vss 0.00857327f
c54 51 Vss 0.00150304f
c55 49 Vss 0.00549985f
c56 47 Vss 0.00136862f
c57 43 Vss 0.00161014f
c58 41 Vss 7.26487e-19
c59 40 Vss 0.00177073f
c60 39 Vss 0.00917963f
c61 38 Vss 0.00784728f
c62 25 Vss 0.085695f
c63 19 Vss 0.0340946f
c64 18 Vss 0.0688517f
c65 8 Vss 0.00226556f
c66 6 Vss 0.0830486f
c67 4 Vss 0.00236553f
c68 2 Vss 0.0834535f
r69 56 59 0.349767
r70 55 56 13.3371
r71 51 59 0.306046
r72 51 53 1.82344
r73 50 57 0.494161
r74 49 55 0.652036
r75 49 50 4.37625
r76 47 65 1.16709
r77 45 57 0.128424
r78 45 47 2.16729
r79 41 43 1.82344
r80 39 57 0.494161
r81 39 40 10.1279
r82 38 41 0.655813
r83 37 40 0.652036
r84 37 38 13.3371
r85 25 65 0.238214
r86 23 25 2.04225
r87 20 23 0.0685365
r88 18 23 0.5835
r89 18 19 2.8008
r90 15 19 0.652036
r91 8 53 1.16709
r92 6 20 2.5674
r93 4 43 1.16709
r94 2 15 2.5674
.ends

.subckt PM_G2_OAI21_N1_B 2 4 10 13 18 21 26 31 Vss
c23 31 Vss 0.00366366f
c24 26 Vss 0.00309808f
c25 18 Vss 6.90549e-19
c26 13 Vss 0.0578401f
c27 2 Vss 0.0576308f
r28 23 31 1.16709
r29 21 23 1.95889
r30 18 26 1.16709
r31 18 21 2.87582
r32 13 31 0.50025
r33 10 26 0.50025
r34 4 13 1.80885
r35 2 10 1.80885
.ends

.subckt PM_G2_OAI21_N1_A 2 4 13 18 26 31 36 43 45 Vss
c43 43 Vss 0.0016451f
c44 36 Vss 0.00277103f
c45 31 Vss 0.00697771f
c46 26 Vss 0.00360766f
c47 18 Vss 0.0860562f
c48 13 Vss 6.71834e-20
c49 4 Vss 0.0575023f
c50 2 Vss 0.0840749f
r51 40 45 0.655813
r52 40 43 9.00257
r53 31 43 1.16709
r54 26 36 1.16709
r55 26 45 4.52212
r56 18 31 0.238214
r57 15 18 1.92555
r58 13 36 0.50025
r59 7 15 0.0685365
r60 4 13 1.80885
r61 2 7 2.5674
.ends

.subckt PM_G2_OAI21_N1_Z 2 4 30 33 Vss
c30 30 Vss 0.00127106f
c31 4 Vss 0.00153036f
c32 2 Vss 0.00148239f
r33 33 35 5.62661
r34 30 33 3.54268
r35 4 35 1.16709
r36 2 30 1.16709
.ends

.subckt PM_G2_OAI21_N1_C 2 4 6 13 14 17 24 27 30 Vss
c30 27 Vss 4.95129e-19
c31 24 Vss 0.0812483f
c32 17 Vss 0.147907f
c33 14 Vss 0.0348316f
c34 13 Vss 0.245605f
c35 4 Vss 0.18102f
c36 2 Vss 0.181207f
r37 27 30 0.0833571
r38 23 24 2.04225
r39 20 24 0.0685365
r40 17 27 1.16709
r41 15 23 0.0685365
r42 15 17 2.8008
r43 13 23 0.5835
r44 13 14 8.92755
r45 10 14 0.652036
r46 6 17 3.0342
r47 4 20 5.835
r48 2 10 5.835
.ends

.subckt G2_OAI21_N1  VSS VDD B A Z C
*
* C	C
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI1.X0 N_Z_XI1.X0_D N_VDD_XI1.X0_PGD N_B_XI1.X0_CG N_C_XI1.X0_PGS N_VSS_XI1.X0_S
+ TIGFET_HPNW1
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_A_XI6.X0_PGS N_VDD_XI6.X0_S
+ TIGFET_HPNW1
XI5.X0 N_Z_XI1.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_C_XI5.X0_PGS N_VSS_XI5.X0_S
+ TIGFET_HPNW1
XI7.X0 N_Z_XI6.X0_D N_VSS_XI7.X0_PGD N_C_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW1
*
x_PM_G2_OAI21_N1_VSS N_VSS_XI1.X0_S N_VSS_XI6.X0_PGD N_VSS_XI5.X0_S
+ N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS N_VSS_c_22_p N_VSS_c_44_p N_VSS_c_1_p
+ N_VSS_c_23_p N_VSS_c_9_p N_VSS_c_24_p N_VSS_c_2_p N_VSS_c_3_p N_VSS_c_7_p
+ N_VSS_c_12_p N_VSS_c_10_p N_VSS_c_16_p VSS Vss PM_G2_OAI21_N1_VSS
x_PM_G2_OAI21_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI6.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI7.X0_S N_VDD_c_50_n N_VDD_c_53_n N_VDD_c_54_n N_VDD_c_55_n
+ N_VDD_c_75_p N_VDD_c_57_n N_VDD_c_60_n N_VDD_c_63_n VDD N_VDD_c_72_p Vss
+ PM_G2_OAI21_N1_VDD
x_PM_G2_OAI21_N1_B N_B_XI1.X0_CG N_B_XI6.X0_CG N_B_c_102_n N_B_c_109_p
+ N_B_c_101_n B N_B_c_105_n N_B_c_107_n Vss PM_G2_OAI21_N1_B
x_PM_G2_OAI21_N1_A N_A_XI6.X0_PGS N_A_XI5.X0_CG N_A_c_139_n N_A_c_149_n
+ N_A_c_125_n N_A_c_127_n N_A_c_131_n A N_A_c_137_n Vss PM_G2_OAI21_N1_A
x_PM_G2_OAI21_N1_Z N_Z_XI1.X0_D N_Z_XI6.X0_D N_Z_c_171_n Z Vss PM_G2_OAI21_N1_Z
x_PM_G2_OAI21_N1_C N_C_XI1.X0_PGS N_C_XI5.X0_PGS N_C_XI7.X0_CG N_C_c_197_n
+ N_C_c_219_n N_C_c_199_n N_C_c_202_n N_C_c_203_n C Vss PM_G2_OAI21_N1_C
cc_1 N_VSS_c_1_p N_VDD_c_50_n 0.00187494f
cc_2 N_VSS_c_2_p N_VDD_c_50_n 0.00510452f
cc_3 N_VSS_c_3_p N_VDD_c_50_n 0.00186257f
cc_4 N_VSS_c_1_p N_VDD_c_53_n 0.0010904f
cc_5 N_VSS_c_2_p N_VDD_c_54_n 0.0014876f
cc_6 N_VSS_c_1_p N_VDD_c_55_n 7.48363e-19
cc_7 N_VSS_c_7_p N_VDD_c_55_n 4.59722e-19
cc_8 N_VSS_XI5.X0_S N_VDD_c_57_n 3.7884e-19
cc_9 N_VSS_c_9_p N_VDD_c_57_n 5.11058e-19
cc_10 N_VSS_c_10_p N_VDD_c_57_n 5.35974e-19
cc_11 N_VSS_c_9_p N_VDD_c_60_n 2.14355e-19
cc_12 N_VSS_c_12_p N_VDD_c_60_n 4.59722e-19
cc_13 N_VSS_c_10_p N_VDD_c_60_n 5.34009e-19
cc_14 N_VSS_c_9_p N_VDD_c_63_n 0.00187494f
cc_15 N_VSS_c_10_p N_VDD_c_63_n 0.00186257f
cc_16 N_VSS_c_16_p N_VDD_c_63_n 0.00730042f
cc_17 N_VSS_c_2_p N_B_c_101_n 5.86846e-19
cc_18 N_VSS_XI6.X0_PGD N_A_XI6.X0_PGS 0.00164631f
cc_19 N_VSS_c_7_p N_A_c_125_n 8.83597e-19
cc_20 N_VSS_c_16_p N_A_c_125_n 4.02032e-19
cc_21 N_VSS_XI6.X0_PGD N_A_c_127_n 3.11814e-19
cc_22 N_VSS_c_22_p N_A_c_127_n 0.00322564f
cc_23 N_VSS_c_23_p N_A_c_127_n 3.44698e-19
cc_24 N_VSS_c_24_p N_A_c_127_n 6.61253e-19
cc_25 N_VSS_c_24_p N_A_c_131_n 3.77503e-19
cc_26 N_VSS_c_23_p A 8.59446e-19
cc_27 N_VSS_c_24_p A 3.44698e-19
cc_28 N_VSS_c_2_p A 0.00272781f
cc_29 N_VSS_c_7_p A 0.00211023f
cc_30 N_VSS_c_16_p A 0.00133784f
cc_31 N_VSS_c_2_p N_A_c_137_n 0.00291082f
cc_32 N_VSS_XI1.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_33 N_VSS_XI5.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_34 N_VSS_c_1_p N_Z_XI1.X0_D 3.48267e-19
cc_35 N_VSS_c_9_p N_Z_XI1.X0_D 3.48267e-19
cc_36 N_VSS_XI1.X0_S N_Z_c_171_n 3.48267e-19
cc_37 N_VSS_XI5.X0_S N_Z_c_171_n 3.48267e-19
cc_38 N_VSS_c_1_p N_Z_c_171_n 5.69026e-19
cc_39 N_VSS_c_9_p N_Z_c_171_n 5.69026e-19
cc_40 N_VSS_c_7_p N_Z_c_171_n 4.84633e-19
cc_41 N_VSS_c_16_p N_Z_c_171_n 4.50981e-19
cc_42 N_VSS_XI6.X0_PGD N_C_c_197_n 6.77138e-19
cc_43 N_VSS_XI7.X0_PGD N_C_c_197_n 6.77138e-19
cc_44 N_VSS_c_44_p N_C_c_199_n 8.9608e-19
cc_45 N_VSS_c_23_p N_C_c_199_n 4.56568e-19
cc_46 N_VSS_c_24_p N_C_c_199_n 0.00315719f
cc_47 N_VSS_XI7.X0_PGS N_C_c_202_n 7.91098e-19
cc_48 N_VSS_c_23_p N_C_c_203_n 5.37794e-19
cc_49 N_VSS_c_24_p N_C_c_203_n 4.56568e-19
cc_50 N_VDD_c_53_n N_B_c_102_n 2.44914e-19
cc_51 N_VDD_c_50_n N_B_c_101_n 0.00216638f
cc_52 N_VDD_c_53_n N_B_c_101_n 2.85486e-19
cc_53 N_VDD_c_50_n N_B_c_105_n 3.66936e-19
cc_54 N_VDD_c_53_n N_B_c_105_n 2.29043e-19
cc_55 N_VDD_c_50_n N_B_c_107_n 4.1997e-19
cc_56 N_VDD_c_72_p N_A_XI5.X0_CG 0.00237871f
cc_57 N_VDD_c_72_p N_A_c_139_n 0.00106215f
cc_58 N_VDD_c_53_n N_A_c_125_n 9.72202e-19
cc_59 N_VDD_c_75_p N_A_c_125_n 7.80108e-19
cc_60 N_VDD_c_63_n N_A_c_125_n 6.23587e-19
cc_61 N_VDD_c_72_p N_A_c_125_n 4.87728e-19
cc_62 N_VDD_c_75_p N_A_c_131_n 4.85469e-19
cc_63 N_VDD_c_63_n N_A_c_131_n 3.66936e-19
cc_64 N_VDD_c_72_p N_A_c_131_n 0.0014909f
cc_65 N_VDD_c_50_n N_A_c_137_n 6.23756e-19
cc_66 N_VDD_c_53_n N_A_c_137_n 2.0345e-19
cc_67 N_VDD_c_53_n N_Z_XI1.X0_D 3.7884e-19
cc_68 N_VDD_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_69 N_VDD_XI7.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_70 N_VDD_c_55_n N_Z_XI6.X0_D 3.72199e-19
cc_71 N_VDD_c_60_n N_Z_XI6.X0_D 3.72199e-19
cc_72 N_VDD_XI6.X0_S N_Z_c_171_n 3.48267e-19
cc_73 N_VDD_XI7.X0_S N_Z_c_171_n 3.48267e-19
cc_74 N_VDD_c_50_n N_Z_c_171_n 3.87755e-19
cc_75 N_VDD_c_53_n N_Z_c_171_n 6.81554e-19
cc_76 N_VDD_c_55_n N_Z_c_171_n 5.6271e-19
cc_77 N_VDD_c_60_n N_Z_c_171_n 7.76033e-19
cc_78 N_VDD_c_63_n N_Z_c_171_n 0.0010014f
cc_79 N_VDD_c_50_n N_C_XI1.X0_PGS 6.09123e-19
cc_80 N_VDD_c_63_n N_C_XI5.X0_PGS 6.28572e-19
cc_81 N_VDD_XI1.X0_PGD N_C_c_197_n 6.72196e-19
cc_82 N_VDD_XI5.X0_PGD N_C_c_197_n 6.76891e-19
cc_83 N_VDD_c_63_n N_C_c_199_n 4.79801e-19
cc_84 N_VDD_c_63_n N_C_c_203_n 3.46645e-19
cc_85 N_B_c_107_n N_A_c_149_n 8.43061e-19
cc_86 N_B_c_109_p N_A_c_127_n 0.00234241f
cc_87 N_B_c_101_n N_A_c_127_n 5.28799e-19
cc_88 N_B_c_107_n N_A_c_127_n 0.00173494f
cc_89 N_B_c_105_n N_A_c_131_n 8.86454e-19
cc_90 N_B_c_101_n A 0.00306515f
cc_91 N_B_c_107_n A 4.56568e-19
cc_92 N_B_c_101_n N_A_c_137_n 6.59436e-19
cc_93 N_B_c_101_n N_Z_c_171_n 0.00673203f
cc_94 N_B_c_105_n N_Z_c_171_n 9.17696e-19
cc_95 N_B_c_107_n N_Z_c_171_n 9.18163e-19
cc_96 N_B_XI1.X0_CG N_C_XI1.X0_PGS 4.42555e-19
cc_97 N_B_c_105_n N_C_XI1.X0_PGS 0.001089f
cc_98 N_B_c_105_n N_C_c_197_n 6.02551e-19
cc_99 N_B_c_107_n N_C_c_197_n 0.00107456f
cc_100 N_B_c_107_n N_C_c_199_n 9.3196e-19
cc_101 N_A_c_125_n N_Z_c_171_n 0.00382179f
cc_102 A N_Z_c_171_n 0.00134325f
cc_103 N_A_XI5.X0_CG N_C_XI5.X0_PGS 4.42555e-19
cc_104 N_A_c_131_n N_C_XI5.X0_PGS 0.001089f
cc_105 N_A_c_131_n N_C_c_197_n 6.59241e-19
cc_106 N_A_XI6.X0_PGS N_C_c_219_n 7.91098e-19
cc_107 N_A_c_125_n N_C_c_199_n 5.38228e-19
cc_108 N_A_c_127_n N_C_c_199_n 2.62413e-19
cc_109 N_A_c_131_n N_C_c_199_n 0.0021499f
cc_110 N_A_c_125_n N_C_c_203_n 8.10255e-19
cc_111 N_Z_c_171_n N_C_c_197_n 4.9701e-19
cc_112 N_Z_c_171_n N_C_c_199_n 9.61365e-19
cc_113 N_Z_c_171_n N_C_c_203_n 0.00143964f
*
.ends
*
*
.subckt OAI21_HPNW1 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 A0 Y B0) G2_OAI21_N1
.ends
*
* File: G3_OR2_N1.pex.netlist
* Created: Tue Mar  1 11:26:38 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_OR2_N1_VSS 2 4 6 10 12 28 29 36 38 52 57 62 67 76 85 90 91 95 96
+ 101 107 113 115 Vss
c75 115 Vss 3.87529e-19
c76 113 Vss 3.75522e-19
c77 107 Vss 0.00356169f
c78 101 Vss 0.00288979f
c79 96 Vss 8.28047e-19
c80 95 Vss 0.00177669f
c81 91 Vss 6.45375e-19
c82 90 Vss 0.00387778f
c83 85 Vss 0.00483971f
c84 76 Vss 0.00487294f
c85 67 Vss 9.52891e-19
c86 62 Vss 6.68032e-19
c87 57 Vss 8.26459e-19
c88 52 Vss 0.00114656f
c89 38 Vss 0.0883089f
c90 36 Vss 6.95992e-20
c91 29 Vss 0.0339709f
c92 28 Vss 0.0988304f
c93 12 Vss 0.0842992f
c94 10 Vss 0.0825208f
c95 6 Vss 0.00148239f
c96 4 Vss 0.0834348f
c97 2 Vss 0.00226843f
r98 108 115 0.494161
r99 107 109 0.652036
r100 107 108 7.46046
r101 103 115 0.128424
r102 102 113 0.494161
r103 101 115 0.494161
r104 101 102 7.46046
r105 97 113 0.128424
r106 95 113 0.494161
r107 95 96 4.37625
r108 90 96 0.652036
r109 89 91 0.655813
r110 89 90 13.3371
r111 67 85 1.16709
r112 67 109 2.16729
r113 62 103 4.83471
r114 57 76 1.16709
r115 57 97 2.16729
r116 52 91 1.82344
r117 36 76 0.238214
r118 36 38 2.04225
r119 31 85 0.238214
r120 29 31 1.45875
r121 28 32 0.652036
r122 28 31 1.45875
r123 25 29 0.652036
r124 22 38 0.0685365
r125 12 32 2.5674
r126 10 25 2.5674
r127 6 62 1.16709
r128 4 22 2.5674
r129 2 52 1.16709
.ends

.subckt PM_G3_OR2_N1_VDD 2 4 6 8 10 12 14 16 37 39 46 49 70 72 73 77 79 83 87 89
+ 93 95 97 102 103 105 106 107 113 119 124 Vss
c84 124 Vss 0.00429743f
c85 119 Vss 0.00559477f
c86 113 Vss 0.00492664f
c87 107 Vss 2.39889e-19
c88 106 Vss 2.39889e-19
c89 103 Vss 3.56526e-19
c90 102 Vss 0.00314642f
c91 97 Vss 0.00307382f
c92 95 Vss 0.00838282f
c93 93 Vss 5.19372e-19
c94 89 Vss 0.00212525f
c95 87 Vss 4.89903e-19
c96 83 Vss 0.00134401f
c97 79 Vss 0.00561519f
c98 77 Vss 0.0016605f
c99 74 Vss 0.00173366f
c100 73 Vss 0.0048947f
c101 72 Vss 0.00279823f
c102 70 Vss 0.00738679f
c103 57 Vss 0.126882f
c104 47 Vss 0.0348458f
c105 46 Vss 0.1003f
c106 39 Vss 7.35265e-20
c107 37 Vss 0.0346129f
c108 36 Vss 0.100535f
c109 16 Vss 0.00262047f
c110 14 Vss 0.0828904f
c111 12 Vss 0.0825208f
c112 10 Vss 0.0828869f
c113 8 Vss 0.0823812f
c114 6 Vss 0.00220666f
c115 4 Vss 0.0830779f
c116 2 Vss 0.0842392f
r117 113 116 0.05
r118 101 102 4.16786
r119 97 101 0.655813
r120 97 99 1.82344
r121 96 107 0.494161
r122 95 102 0.652036
r123 95 96 10.1279
r124 93 124 1.16709
r125 91 107 0.128424
r126 91 93 2.16729
r127 90 106 0.494161
r128 89 107 0.494161
r129 89 90 4.54296
r130 87 119 1.16709
r131 85 106 0.128424
r132 85 87 2.16729
r133 83 116 1.16709
r134 81 83 2.20896
r135 80 105 0.326018
r136 79 106 0.494161
r137 79 80 10.1696
r138 75 103 0.0828784
r139 75 77 1.82344
r140 73 81 0.652036
r141 73 74 4.37625
r142 72 105 0.326018
r143 71 103 0.551426
r144 71 72 4.16786
r145 70 103 0.551426
r146 69 74 0.652036
r147 69 70 13.3371
r148 56 113 0.262036
r149 56 57 2.26917
r150 53 56 2.26917
r151 49 124 0.238214
r152 47 49 1.45875
r153 46 50 0.652036
r154 46 49 1.45875
r155 43 47 0.652036
r156 39 119 0.238214
r157 37 39 1.5171
r158 36 40 0.652036
r159 36 39 1.4004
r160 33 37 0.652036
r161 30 57 0.00605528
r162 27 53 0.00605528
r163 16 99 1.16709
r164 14 43 2.5674
r165 12 50 2.5674
r166 10 40 2.5674
r167 8 33 2.5674
r168 6 77 1.16709
r169 4 27 2.5674
r170 2 30 2.5674
.ends

.subckt PM_G3_OR2_N1_B 2 4 10 13 18 21 26 31 Vss
c25 31 Vss 0.00183593f
c26 26 Vss 0.00362926f
c27 18 Vss 0.00110935f
c28 13 Vss 0.057478f
c29 10 Vss 6.71834e-20
c30 2 Vss 0.0576626f
r31 23 31 1.16709
r32 21 23 2.08393
r33 18 26 1.16709
r34 18 21 2.75079
r35 13 31 0.50025
r36 10 26 0.50025
r37 4 13 1.80885
r38 2 10 1.80885
.ends

.subckt PM_G3_OR2_N1_NET21 2 4 8 10 21 24 45 53 66 70 Vss
c39 70 Vss 0.00761723f
c40 66 Vss 0.00611981f
c41 53 Vss 0.00155023f
c42 45 Vss 0.00245986f
c43 24 Vss 0.225594f
c44 21 Vss 0.0713786f
c45 19 Vss 0.0247918f
c46 10 Vss 0.0847975f
c47 4 Vss 0.00148239f
c48 2 Vss 0.0021264f
r49 70 74 0.652036
r50 53 66 1.16709
r51 53 74 2.9175
r52 48 70 8.04396
r53 48 50 5.66829
r54 45 48 3.501
r55 27 66 0.0476429
r56 25 27 0.326018
r57 25 27 0.1167
r58 24 28 0.652036
r59 24 27 6.7686
r60 21 66 0.357321
r61 19 27 0.326018
r62 19 21 0.40845
r63 10 28 2.5674
r64 8 21 2.15895
r65 4 50 1.16709
r66 2 45 1.16709
.ends

.subckt PM_G3_OR2_N1_A 2 4 10 11 14 18 Vss
c22 18 Vss 2.95942e-19
c23 14 Vss 0.116245f
c24 11 Vss 0.0348164f
c25 10 Vss 0.273261f
c26 2 Vss 0.142908f
r27 21 27 1.16709
r28 18 21 0.0833571
r29 14 27 0.05
r30 12 14 1.6338
r31 10 12 0.652036
r32 10 11 8.92755
r33 7 11 0.652036
r34 4 14 3.0342
r35 2 7 4.668
.ends

.subckt PM_G3_OR2_N1_Z 2 16 19 Vss
c11 2 Vss 0.00148239f
r12 16 19 0.0364688
r13 2 19 1.16709
.ends

.subckt G3_OR2_N1  VSS VDD B A Z
*
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI2.X0 N_NET21_XI2.X0_D N_VDD_XI2.X0_PGD N_B_XI2.X0_CG N_VDD_XI2.X0_PGS
+ N_VSS_XI2.X0_S TIGFET_HPNW1
XI0.X0 N_NET21_XI0.X0_D N_VSS_XI0.X0_PGD N_B_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW1
XI1.X0 N_NET21_XI0.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_NET21_XI3.X0_CG N_VDD_XI3.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW1
XI4.X0 N_Z_XI3.X0_D N_VSS_XI4.X0_PGD N_NET21_XI4.X0_CG N_VSS_XI4.X0_PGS
+ N_VDD_XI4.X0_S TIGFET_HPNW1
*
x_PM_G3_OR2_N1_VSS N_VSS_XI2.X0_S N_VSS_XI0.X0_PGD N_VSS_XI1.X0_S
+ N_VSS_XI4.X0_PGD N_VSS_XI4.X0_PGS N_VSS_c_32_p N_VSS_c_4_p N_VSS_c_51_p
+ N_VSS_c_3_p N_VSS_c_6_p N_VSS_c_9_p N_VSS_c_23_p N_VSS_c_30_p N_VSS_c_10_p
+ N_VSS_c_31_p N_VSS_c_7_p N_VSS_c_8_p N_VSS_c_19_p N_VSS_c_12_p N_VSS_c_20_p
+ N_VSS_c_27_p N_VSS_c_21_p VSS Vss PM_G3_OR2_N1_VSS
x_PM_G3_OR2_N1_VDD N_VDD_XI2.X0_PGD N_VDD_XI2.X0_PGS N_VDD_XI0.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI3.X0_PGD N_VDD_XI3.X0_PGS
+ N_VDD_XI4.X0_S N_VDD_c_78_n N_VDD_c_149_p N_VDD_c_79_n N_VDD_c_140_p
+ N_VDD_c_80_n N_VDD_c_84_n N_VDD_c_88_n N_VDD_c_90_n N_VDD_c_91_n N_VDD_c_124_p
+ N_VDD_c_97_n N_VDD_c_100_n N_VDD_c_104_n N_VDD_c_107_n N_VDD_c_156_p
+ N_VDD_c_112_n N_VDD_c_114_n VDD N_VDD_c_115_n N_VDD_c_116_n N_VDD_c_121_p
+ N_VDD_c_117_n N_VDD_c_119_n Vss PM_G3_OR2_N1_VDD
x_PM_G3_OR2_N1_B N_B_XI2.X0_CG N_B_XI0.X0_CG N_B_c_169_n N_B_c_160_n N_B_c_161_n
+ B N_B_c_164_n N_B_c_165_n Vss PM_G3_OR2_N1_B
x_PM_G3_OR2_N1_NET21 N_NET21_XI2.X0_D N_NET21_XI0.X0_D N_NET21_XI3.X0_CG
+ N_NET21_XI4.X0_CG N_NET21_c_203_n N_NET21_c_190_n N_NET21_c_191_n
+ N_NET21_c_195_n N_NET21_c_212_n N_NET21_c_197_n Vss PM_G3_OR2_N1_NET21
x_PM_G3_OR2_N1_A N_A_XI0.X0_PGS N_A_XI1.X0_CG N_A_c_224_n N_A_c_228_n
+ N_A_c_230_n A Vss PM_G3_OR2_N1_A
x_PM_G3_OR2_N1_Z N_Z_XI3.X0_D Z N_Z_c_248_n Vss PM_G3_OR2_N1_Z
cc_1 N_VSS_XI0.X0_PGD N_VDD_XI1.X0_PGD 0.00175996f
cc_2 N_VSS_XI4.X0_PGD N_VDD_XI3.X0_PGD 0.00168578f
cc_3 N_VSS_c_3_p N_VDD_c_78_n 0.00175996f
cc_4 N_VSS_c_4_p N_VDD_c_79_n 0.00168578f
cc_5 N_VSS_XI2.X0_S N_VDD_c_80_n 9.5668e-19
cc_6 N_VSS_c_6_p N_VDD_c_80_n 0.00165395f
cc_7 N_VSS_c_7_p N_VDD_c_80_n 0.00519974f
cc_8 N_VSS_c_8_p N_VDD_c_80_n 0.00186257f
cc_9 N_VSS_c_9_p N_VDD_c_84_n 4.43871e-19
cc_10 N_VSS_c_10_p N_VDD_c_84_n 3.66936e-19
cc_11 N_VSS_c_7_p N_VDD_c_84_n 0.00303537f
cc_12 N_VSS_c_12_p N_VDD_c_84_n 0.00106607f
cc_13 N_VSS_XI2.X0_S N_VDD_c_88_n 3.7884e-19
cc_14 N_VSS_c_6_p N_VDD_c_88_n 0.00104703f
cc_15 N_VSS_c_6_p N_VDD_c_90_n 7.47067e-19
cc_16 N_VSS_c_3_p N_VDD_c_91_n 3.37151e-19
cc_17 N_VSS_c_9_p N_VDD_c_91_n 0.00161703f
cc_18 N_VSS_c_10_p N_VDD_c_91_n 2.03837e-19
cc_19 N_VSS_c_19_p N_VDD_c_91_n 0.0034844f
cc_20 N_VSS_c_20_p N_VDD_c_91_n 0.00432568f
cc_21 N_VSS_c_21_p N_VDD_c_91_n 7.74609e-19
cc_22 N_VSS_c_9_p N_VDD_c_97_n 8.45115e-19
cc_23 N_VSS_c_23_p N_VDD_c_97_n 3.93845e-19
cc_24 N_VSS_c_10_p N_VDD_c_97_n 3.95933e-19
cc_25 N_VSS_c_23_p N_VDD_c_100_n 5.01863e-19
cc_26 N_VSS_c_20_p N_VDD_c_100_n 0.00137553f
cc_27 N_VSS_c_27_p N_VDD_c_100_n 0.00142235f
cc_28 VSS N_VDD_c_100_n 0.00104966f
cc_29 N_VSS_c_23_p N_VDD_c_104_n 3.91951e-19
cc_30 N_VSS_c_30_p N_VDD_c_104_n 8.51944e-19
cc_31 N_VSS_c_31_p N_VDD_c_104_n 3.99794e-19
cc_32 N_VSS_c_32_p N_VDD_c_107_n 3.80388e-19
cc_33 N_VSS_c_4_p N_VDD_c_107_n 3.60588e-19
cc_34 N_VSS_c_30_p N_VDD_c_107_n 0.00141604f
cc_35 N_VSS_c_31_p N_VDD_c_107_n 0.00112293f
cc_36 N_VSS_c_27_p N_VDD_c_107_n 0.00608608f
cc_37 N_VSS_c_30_p N_VDD_c_112_n 9.12964e-19
cc_38 N_VSS_c_31_p N_VDD_c_112_n 3.66936e-19
cc_39 N_VSS_c_7_p N_VDD_c_114_n 0.00116512f
cc_40 N_VSS_c_20_p N_VDD_c_115_n 9.75006e-19
cc_41 N_VSS_c_27_p N_VDD_c_116_n 9.68945e-19
cc_42 N_VSS_c_9_p N_VDD_c_117_n 3.44698e-19
cc_43 N_VSS_c_10_p N_VDD_c_117_n 7.93802e-19
cc_44 N_VSS_c_30_p N_VDD_c_119_n 3.48267e-19
cc_45 N_VSS_c_31_p N_VDD_c_119_n 8.07896e-19
cc_46 N_VSS_c_10_p N_B_c_160_n 0.00234321f
cc_47 N_VSS_c_9_p N_B_c_161_n 8.39582e-19
cc_48 N_VSS_c_10_p N_B_c_161_n 5.42695e-19
cc_49 N_VSS_c_7_p N_B_c_161_n 7.94601e-19
cc_50 N_VSS_c_10_p N_B_c_164_n 2.00604e-19
cc_51 N_VSS_c_51_p N_B_c_165_n 8.37306e-19
cc_52 N_VSS_c_9_p N_B_c_165_n 4.56568e-19
cc_53 N_VSS_c_10_p N_B_c_165_n 0.00173573f
cc_54 N_VSS_XI2.X0_S N_NET21_XI2.X0_D 3.43419e-19
cc_55 N_VSS_c_6_p N_NET21_XI2.X0_D 3.48267e-19
cc_56 N_VSS_XI1.X0_S N_NET21_XI0.X0_D 3.43419e-19
cc_57 N_VSS_c_23_p N_NET21_XI0.X0_D 3.48267e-19
cc_58 N_VSS_c_31_p N_NET21_XI4.X0_CG 7.99056e-19
cc_59 N_VSS_XI4.X0_PGD N_NET21_c_190_n 4.20799e-19
cc_60 N_VSS_XI1.X0_S N_NET21_c_191_n 3.48267e-19
cc_61 N_VSS_c_6_p N_NET21_c_191_n 8.89782e-19
cc_62 N_VSS_c_23_p N_NET21_c_191_n 5.69026e-19
cc_63 N_VSS_c_7_p N_NET21_c_191_n 2.81358e-19
cc_64 N_VSS_c_7_p N_NET21_c_195_n 2.56803e-19
cc_65 N_VSS_c_27_p N_NET21_c_195_n 2.99166e-19
cc_66 N_VSS_c_23_p N_NET21_c_197_n 9.55513e-19
cc_67 N_VSS_c_7_p N_NET21_c_197_n 2.03357e-19
cc_68 N_VSS_c_20_p N_NET21_c_197_n 9.1856e-19
cc_69 N_VSS_XI0.X0_PGD N_A_c_224_n 9.39677e-19
cc_70 N_VSS_c_3_p N_A_c_224_n 2.16729e-19
cc_71 N_VSS_XI1.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_72 N_VSS_c_23_p N_Z_XI3.X0_D 3.48267e-19
cc_73 N_VSS_XI1.X0_S N_Z_c_248_n 3.48267e-19
cc_74 N_VSS_c_23_p N_Z_c_248_n 7.85754e-19
cc_75 N_VSS_c_27_p N_Z_c_248_n 2.64173e-19
cc_76 N_VDD_c_121_p N_B_XI2.X0_CG 0.00237871f
cc_77 N_VDD_c_121_p N_B_c_169_n 0.00105622f
cc_78 N_VDD_c_80_n N_B_c_161_n 0.0025613f
cc_79 N_VDD_c_124_p N_B_c_161_n 7.31965e-19
cc_80 N_VDD_c_121_p N_B_c_161_n 5.48584e-19
cc_81 N_VDD_c_80_n N_B_c_164_n 4.9897e-19
cc_82 N_VDD_c_124_p N_B_c_164_n 4.85469e-19
cc_83 N_VDD_c_121_p N_B_c_164_n 0.00150793f
cc_84 N_VDD_c_80_n N_B_c_165_n 3.66936e-19
cc_85 N_VDD_c_121_p N_B_c_165_n 2.00604e-19
cc_86 N_VDD_XI0.X0_S N_NET21_XI0.X0_D 3.43419e-19
cc_87 N_VDD_c_90_n N_NET21_XI0.X0_D 3.72199e-19
cc_88 N_VDD_c_91_n N_NET21_XI0.X0_D 3.7884e-19
cc_89 N_VDD_c_119_n N_NET21_c_203_n 0.00250475f
cc_90 N_VDD_XI3.X0_PGD N_NET21_c_190_n 4.25379e-19
cc_91 N_VDD_XI0.X0_S N_NET21_c_191_n 3.48267e-19
cc_92 N_VDD_c_80_n N_NET21_c_191_n 4.38672e-19
cc_93 N_VDD_c_90_n N_NET21_c_191_n 7.89245e-19
cc_94 N_VDD_c_91_n N_NET21_c_191_n 5.36364e-19
cc_95 N_VDD_c_140_p N_NET21_c_195_n 3.64358e-19
cc_96 N_VDD_c_104_n N_NET21_c_195_n 6.84156e-19
cc_97 N_VDD_c_119_n N_NET21_c_195_n 4.99367e-19
cc_98 N_VDD_c_104_n N_NET21_c_212_n 4.85469e-19
cc_99 N_VDD_c_119_n N_NET21_c_212_n 0.0014909f
cc_100 N_VDD_XI2.X0_PGD N_A_c_224_n 5.10213e-19
cc_101 N_VDD_XI1.X0_PGD N_A_c_224_n 2.48727e-19
cc_102 N_VDD_XI2.X0_PGS N_A_c_228_n 6.4837e-19
cc_103 N_VDD_c_80_n N_A_c_228_n 3.16598e-19
cc_104 N_VDD_c_149_p N_A_c_230_n 8.9931e-19
cc_105 N_VDD_c_97_n N_A_c_230_n 4.91217e-19
cc_106 N_VDD_c_117_n N_A_c_230_n 0.00142365f
cc_107 N_VDD_c_97_n A 6.02732e-19
cc_108 N_VDD_c_117_n A 4.56568e-19
cc_109 N_VDD_XI4.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_110 N_VDD_c_107_n N_Z_XI3.X0_D 3.7884e-19
cc_111 N_VDD_c_156_p N_Z_XI3.X0_D 3.72199e-19
cc_112 N_VDD_XI4.X0_S N_Z_c_248_n 3.48267e-19
cc_113 N_VDD_c_107_n N_Z_c_248_n 5.12447e-19
cc_114 N_VDD_c_156_p N_Z_c_248_n 7.4527e-19
cc_115 N_B_c_161_n N_NET21_c_191_n 0.00757794f
cc_116 N_B_c_164_n N_NET21_c_191_n 9.56873e-19
cc_117 N_B_c_165_n N_NET21_c_191_n 8.92526e-19
cc_118 N_B_c_160_n N_A_XI0.X0_PGS 4.5346e-19
cc_119 N_B_c_165_n N_A_XI0.X0_PGS 7.86826e-19
cc_120 N_B_c_164_n N_A_c_224_n 9.25308e-19
cc_121 N_B_c_165_n N_A_c_230_n 7.50183e-19
cc_122 N_NET21_c_191_n N_A_c_224_n 8.63036e-19
cc_123 N_NET21_c_191_n N_A_c_230_n 9.38449e-19
cc_124 N_NET21_c_195_n N_A_c_230_n 3.48267e-19
cc_125 N_NET21_c_212_n N_A_c_230_n 0.00196751f
cc_126 N_NET21_c_191_n A 0.00142917f
cc_127 N_NET21_c_195_n A 4.28721e-19
cc_128 N_NET21_c_197_n A 3.26205e-19
*
.ends
*
*
.subckt OR2_HPNW1 A B Y VDD VSS
xgate (VSS VDD B A Y) G3_OR2_N1
.ends
*
* File: G4_XNOR2_N1.pex.netlist
* Created: Wed Mar 16 10:29:55 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XNOR2_N1_VDD 2 5 9 12 16 32 35 42 43 66 68 69 70 73 75 76 79 81 85
+ 89 91 93 98 99 100 103 109 114 Vss
c113 114 Vss 0.00462632f
c114 109 Vss 0.00491723f
c115 101 Vss 8.54719e-19
c116 100 Vss 2.39889e-19
c117 99 Vss 3.56526e-19
c118 98 Vss 0.0049606f
c119 93 Vss 0.00247173f
c120 91 Vss 0.0107823f
c121 89 Vss 0.00155915f
c122 85 Vss 3.94646e-19
c123 81 Vss 0.00431979f
c124 79 Vss 0.00104496f
c125 76 Vss 8.67334e-19
c126 75 Vss 0.00219831f
c127 73 Vss 0.00159894f
c128 70 Vss 8.63261e-19
c129 69 Vss 0.00531705f
c130 68 Vss 0.00645016f
c131 66 Vss 0.00203422f
c132 43 Vss 0.0336444f
c133 42 Vss 0.0994765f
c134 35 Vss 7.78608e-20
c135 33 Vss 0.0348624f
c136 32 Vss 0.0999592f
c137 16 Vss 0.00272748f
c138 12 Vss 0.00264503f
c139 9 Vss 0.165252f
c140 5 Vss 0.165777f
c141 2 Vss 0.00272748f
r142 98 103 0.326018
r143 97 98 4.16786
r144 93 97 0.655813
r145 93 95 1.82344
r146 92 101 0.494161
r147 91 103 0.326018
r148 91 92 13.0037
r149 87 101 0.128424
r150 87 89 4.83471
r151 85 114 1.16709
r152 83 85 2.16729
r153 82 100 0.494161
r154 81 101 0.494161
r155 81 82 7.46046
r156 79 109 1.16709
r157 77 100 0.128424
r158 77 79 2.16729
r159 75 100 0.494161
r160 75 76 4.37625
r161 71 99 0.0828784
r162 71 73 1.82344
r163 69 83 0.652036
r164 69 70 10.1279
r165 68 76 0.652036
r166 67 99 0.551426
r167 67 68 12.1701
r168 66 99 0.551426
r169 65 70 0.652036
r170 65 66 4.16786
r171 45 114 0.238214
r172 43 45 1.45875
r173 42 46 0.652036
r174 42 45 1.45875
r175 39 43 0.652036
r176 35 109 0.238214
r177 33 35 1.45875
r178 32 36 0.652036
r179 32 35 1.45875
r180 29 33 0.652036
r181 16 95 1.16709
r182 12 89 1.16709
r183 9 46 2.5674
r184 9 39 2.5674
r185 5 36 2.5674
r186 5 29 2.5674
r187 2 73 1.16709
.ends

.subckt PM_G4_XNOR2_N1_VSS 3 6 8 11 16 32 33 42 43 66 71 76 81 87 96 101 114 116
+ 117 118 123 124 129 137 142 143 144 146 Vss
c99 144 Vss 3.75522e-19
c100 143 Vss 3.21033e-19
c101 142 Vss 0.00224529f
c102 141 Vss 0.0013489f
c103 137 Vss 0.00215359f
c104 129 Vss 0.0112621f
c105 124 Vss 8.17415e-19
c106 123 Vss 0.00403195f
c107 118 Vss 8.39382e-19
c108 117 Vss 0.00163605f
c109 116 Vss 0.00144702f
c110 114 Vss 0.00415033f
c111 101 Vss 0.00449981f
c112 96 Vss 0.00516182f
c113 87 Vss 7.10513e-22
c114 81 Vss 0.00255515f
c115 76 Vss 9.53239e-19
c116 71 Vss 0.00133653f
c117 66 Vss 0.00143917f
c118 43 Vss 0.033325f
c119 42 Vss 0.0990666f
c120 33 Vss 0.0336725f
c121 32 Vss 0.0976281f
c122 16 Vss 0.00213567f
c123 11 Vss 0.165384f
c124 8 Vss 0.00163738f
c125 6 Vss 0.00213969f
c126 3 Vss 0.166856f
r127 141 146 0.326018
r128 141 142 4.16786
r129 137 142 0.655813
r130 130 144 0.494161
r131 129 146 0.326018
r132 125 144 0.128424
r133 123 133 0.652036
r134 123 124 10.1279
r135 119 143 0.0828784
r136 117 144 0.494161
r137 117 118 4.37625
r138 116 124 0.652036
r139 115 143 0.551426
r140 115 116 4.16786
r141 114 143 0.551426
r142 113 118 0.652036
r143 113 114 12.1701
r144 87 137 1.82344
r145 81 129 13.5872
r146 81 130 8.04396
r147 81 84 5.37654
r148 76 101 1.16709
r149 76 133 2.16729
r150 71 96 1.16709
r151 71 125 2.16729
r152 66 119 1.82344
r153 45 101 0.238214
r154 43 45 1.45875
r155 42 46 0.652036
r156 42 45 1.45875
r157 39 43 0.652036
r158 35 96 0.238214
r159 33 35 1.45875
r160 32 36 0.652036
r161 32 35 1.45875
r162 29 33 0.652036
r163 16 87 1.16709
r164 11 46 2.5674
r165 11 39 2.5674
r166 8 84 1.16709
r167 6 66 1.16709
r168 3 36 2.5674
r169 3 29 2.5674
.ends

.subckt PM_G4_XNOR2_N1_A 2 4 7 10 18 21 24 28 39 48 51 54 57 62 67 72 77 85 Vss
c60 85 Vss 9.00557e-19
c61 77 Vss 0.00241581f
c62 72 Vss 0.00594049f
c63 67 Vss 0.00360869f
c64 62 Vss 0.00199403f
c65 57 Vss 0.00406361f
c66 51 Vss 8.38354e-19
c67 48 Vss 0.124108f
c68 43 Vss 0.0295947f
c69 39 Vss 4.97883e-20
c70 28 Vss 0.152592f
c71 24 Vss 2.44824e-19
c72 21 Vss 0.169386f
c73 18 Vss 0.0714048f
c74 16 Vss 0.0247918f
c75 10 Vss 0.0674191f
c76 7 Vss 0.219196f
c77 4 Vss 0.08397f
r78 81 85 0.653045
r79 62 77 1.16709
r80 62 85 4.9014
r81 57 72 1.16709
r82 57 81 7.87725
r83 51 67 1.16709
r84 51 54 0.0416786
r85 47 72 0.262036
r86 47 48 2.334
r87 44 47 2.20433
r88 39 77 0.404964
r89 33 48 0.00605528
r90 31 44 0.00605528
r91 29 43 0.494161
r92 28 30 0.652036
r93 28 29 4.84305
r94 25 43 0.128424
r95 24 67 0.0476429
r96 22 24 0.326018
r97 22 24 0.1167
r98 21 43 0.494161
r99 21 24 6.7686
r100 18 67 0.357321
r101 16 24 0.326018
r102 16 18 0.40845
r103 10 39 2.04225
r104 7 33 2.5674
r105 7 31 2.5674
r106 7 30 2.5674
r107 4 25 2.5674
r108 2 18 2.15895
.ends

.subckt PM_G4_XNOR2_N1_NET1 2 7 10 31 35 44 49 58 66 Vss
c38 66 Vss 6.40075e-20
c39 58 Vss 0.00598766f
c40 49 Vss 0.00482775f
c41 44 Vss 0.00129308f
c42 35 Vss 0.126399f
c43 31 Vss 0.128923f
c44 10 Vss 0.135805f
c45 7 Vss 0.297098f
c46 2 Vss 0.0015894f
r47 62 66 0.653045
r48 49 58 1.16709
r49 49 66 12.9148
r50 44 62 2.08393
r51 33 35 1.45875
r52 30 58 0.262036
r53 30 31 2.20433
r54 27 30 2.334
r55 25 35 0.259088
r56 24 31 0.00605528
r57 21 33 0.259088
r58 18 27 0.00605528
r59 10 21 4.25955
r60 7 25 5.30985
r61 7 24 2.5674
r62 7 18 2.5674
r63 2 44 1.16709
.ends

.subckt PM_G4_XNOR2_N1_NET2 2 6 9 21 22 33 42 47 56 74 Vss
c50 74 Vss 3.88292e-19
c51 56 Vss 0.00473316f
c52 47 Vss 0.00694068f
c53 42 Vss 0.00195908f
c54 33 Vss 0.123617f
c55 22 Vss 0.0344905f
c56 21 Vss 0.177827f
c57 9 Vss 0.362751f
c58 6 Vss 0.0802803f
c59 2 Vss 0.0015894f
r60 70 74 0.660011
r61 47 56 1.16709
r62 47 74 11.3611
r63 42 70 1.95889
r64 32 56 0.262036
r65 32 33 2.26917
r66 29 32 2.26917
r67 26 33 0.00605528
r68 24 29 0.00605528
r69 21 23 0.652036
r70 21 22 4.84305
r71 18 22 0.652036
r72 9 26 2.5674
r73 9 24 2.5674
r74 9 23 7.4688
r75 6 18 2.5674
r76 2 42 1.16709
.ends

.subckt PM_G4_XNOR2_N1_B 2 4 7 10 19 20 28 33 37 38 48 52 55 58 61 Vss
c37 61 Vss 0.0280185f
c38 55 Vss 9.41292e-19
c39 52 Vss 0.134888f
c40 48 Vss 0.0597924f
c41 38 Vss 0.0333789f
c42 37 Vss 0.090068f
c43 33 Vss 0.0345164f
c44 28 Vss 0.0897381f
c45 20 Vss 0.0343755f
c46 19 Vss 0.169386f
c47 10 Vss 0.155214f
c48 7 Vss 0.216f
c49 4 Vss 0.0714224f
c50 2 Vss 0.0847975f
r51 55 61 1.16709
r52 55 58 0.166714
r53 50 52 4.53833
r54 47 48 1.167
r55 42 52 0.00605528
r56 37 39 0.652036
r57 37 38 2.04225
r58 35 48 0.0685365
r59 34 50 0.00605528
r60 33 38 0.652036
r61 32 47 0.0685365
r62 32 33 1.2837
r63 31 61 0.181909
r64 29 61 0.494161
r65 29 31 0.1167
r66 28 47 0.5835
r67 28 31 3.55935
r68 23 61 0.128424
r69 23 61 0.40845
r70 22 61 0.181909
r71 20 22 6.7686
r72 19 61 0.494161
r73 19 22 0.1167
r74 16 20 0.652036
r75 10 39 5.0181
r76 7 42 2.5674
r77 7 35 2.5674
r78 7 34 2.5674
r79 4 61 2.15895
r80 2 16 2.5674
.ends

.subckt PM_G4_XNOR2_N1_Z 2 4 30 33 Vss
c27 30 Vss 0.00253242f
c28 4 Vss 0.00249005f
c29 2 Vss 0.00153036f
r30 33 35 2.9175
r31 30 33 5.08479
r32 4 35 1.16709
r33 2 30 1.16709
.ends

.subckt G4_XNOR2_N1  VDD VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI1.X0 N_NET1_XI1.X0_D N_VSS_XI1.X0_PGD N_B_XI1.X0_CG N_VSS_XI1.X0_PGD
+ N_VDD_XI1.X0_S TIGFET_HPNW1
XI9.X0 N_NET2_XI9.X0_D N_VDD_XI9.X0_PGD N_A_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW1
XI10.X0 N_NET1_XI1.X0_D N_VDD_XI10.X0_PGD N_B_XI10.X0_CG N_VDD_XI10.X0_PGD
+ N_VSS_XI10.X0_S TIGFET_HPNW1
XI3.X0 N_NET2_XI9.X0_D N_VSS_XI3.X0_PGD N_A_XI3.X0_CG N_VSS_XI3.X0_PGD
+ N_VDD_XI3.X0_S TIGFET_HPNW1
XI5.X0 N_Z_XI5.X0_D N_B_XI5.X0_PGD N_NET2_XI5.X0_CG N_B_XI5.X0_PGD
+ N_VSS_XI10.X0_S TIGFET_HPNW1
XI8.X0 N_Z_XI8.X0_D N_A_XI8.X0_PGD N_B_XI8.X0_CG N_A_XI8.X0_PGD N_VDD_XI3.X0_S
+ TIGFET_HPNW1
XI11.X0 N_Z_XI5.X0_D N_NET1_XI11.X0_PGD N_A_XI11.X0_CG N_NET1_XI11.X0_PGD
+ N_VSS_XI11.X0_S TIGFET_HPNW1
XI7.X0 N_Z_XI8.X0_D N_NET2_XI7.X0_PGD N_NET1_XI7.X0_CG N_NET2_XI7.X0_PGD
+ N_VDD_XI7.X0_S TIGFET_HPNW1
*
x_PM_G4_XNOR2_N1_VDD N_VDD_XI1.X0_S N_VDD_XI9.X0_PGD N_VDD_XI10.X0_PGD
+ N_VDD_XI3.X0_S N_VDD_XI7.X0_S N_VDD_c_11_p N_VDD_c_58_p N_VDD_c_26_p
+ N_VDD_c_8_p N_VDD_c_17_p N_VDD_c_14_p N_VDD_c_9_p N_VDD_c_45_p N_VDD_c_3_p
+ N_VDD_c_16_p N_VDD_c_49_p N_VDD_c_21_p N_VDD_c_12_p N_VDD_c_19_p N_VDD_c_4_p
+ N_VDD_c_60_p N_VDD_c_7_p N_VDD_c_90_p N_VDD_c_42_p N_VDD_c_48_p VDD
+ N_VDD_c_24_p N_VDD_c_20_p Vss PM_G4_XNOR2_N1_VDD
x_PM_G4_XNOR2_N1_VSS N_VSS_XI1.X0_PGD N_VSS_XI9.X0_S N_VSS_XI10.X0_S
+ N_VSS_XI3.X0_PGD N_VSS_XI11.X0_S N_VSS_c_121_n N_VSS_c_123_n N_VSS_c_172_p
+ N_VSS_c_124_n N_VSS_c_126_n N_VSS_c_130_n N_VSS_c_134_n N_VSS_c_138_n
+ N_VSS_c_143_n N_VSS_c_145_n N_VSS_c_149_n N_VSS_c_153_n N_VSS_c_156_n
+ N_VSS_c_157_n N_VSS_c_158_n N_VSS_c_159_n N_VSS_c_162_n N_VSS_c_163_n
+ N_VSS_c_164_n N_VSS_c_185_p N_VSS_c_165_n N_VSS_c_166_n VSS Vss
+ PM_G4_XNOR2_N1_VSS
x_PM_G4_XNOR2_N1_A N_A_XI9.X0_CG N_A_XI3.X0_CG N_A_XI8.X0_PGD N_A_XI11.X0_CG
+ N_A_c_214_n N_A_c_215_n N_A_c_217_n N_A_c_218_n N_A_c_249_p N_A_c_219_n
+ N_A_c_220_n A N_A_c_223_n N_A_c_225_n N_A_c_226_n N_A_c_229_n N_A_c_244_p
+ N_A_c_242_n Vss PM_G4_XNOR2_N1_A
x_PM_G4_XNOR2_N1_NET1 N_NET1_XI1.X0_D N_NET1_XI11.X0_PGD N_NET1_XI7.X0_CG
+ N_NET1_c_309_p N_NET1_c_293_n N_NET1_c_276_n N_NET1_c_279_n N_NET1_c_296_n
+ N_NET1_c_280_n Vss PM_G4_XNOR2_N1_NET1
x_PM_G4_XNOR2_N1_NET2 N_NET2_XI9.X0_D N_NET2_XI5.X0_CG N_NET2_XI7.X0_PGD
+ N_NET2_c_336_n N_NET2_c_356_p N_NET2_c_314_n N_NET2_c_315_n N_NET2_c_318_n
+ N_NET2_c_322_n N_NET2_c_324_n Vss PM_G4_XNOR2_N1_NET2
x_PM_G4_XNOR2_N1_B N_B_XI1.X0_CG N_B_XI10.X0_CG N_B_XI5.X0_PGD N_B_XI8.X0_CG
+ N_B_c_363_n N_B_c_382_n N_B_c_365_n N_B_c_392_n N_B_c_388_n N_B_c_384_n
+ N_B_c_395_n N_B_c_366_n N_B_c_367_n B N_B_c_369_n Vss PM_G4_XNOR2_N1_B
x_PM_G4_XNOR2_N1_Z N_Z_XI5.X0_D N_Z_XI8.X0_D N_Z_c_403_n Z Vss PM_G4_XNOR2_N1_Z
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI1.X0_PGD 2.96813e-19
cc_2 N_VDD_XI10.X0_PGD N_VSS_XI1.X0_PGD 0.00168295f
cc_3 N_VDD_c_3_p N_VSS_XI9.X0_S 2.15082e-19
cc_4 N_VDD_c_4_p N_VSS_XI10.X0_S 2.35318e-19
cc_5 N_VDD_XI9.X0_PGD N_VSS_XI3.X0_PGD 0.00167677f
cc_6 N_VDD_c_4_p N_VSS_XI3.X0_PGD 2.68479e-19
cc_7 N_VDD_c_7_p N_VSS_XI11.X0_S 2.15082e-19
cc_8 N_VDD_c_8_p N_VSS_c_121_n 0.00168295f
cc_9 N_VDD_c_9_p N_VSS_c_121_n 3.60588e-19
cc_10 N_VDD_c_9_p N_VSS_c_123_n 3.60588e-19
cc_11 N_VDD_c_11_p N_VSS_c_124_n 0.00167677f
cc_12 N_VDD_c_12_p N_VSS_c_124_n 3.60588e-19
cc_13 N_VDD_XI1.X0_S N_VSS_c_126_n 2.15082e-19
cc_14 N_VDD_c_14_p N_VSS_c_126_n 0.00187494f
cc_15 N_VDD_c_3_p N_VSS_c_126_n 8.9077e-19
cc_16 N_VDD_c_16_p N_VSS_c_126_n 5.16845e-19
cc_17 N_VDD_c_17_p N_VSS_c_130_n 4.43871e-19
cc_18 N_VDD_c_9_p N_VSS_c_130_n 0.00141228f
cc_19 N_VDD_c_19_p N_VSS_c_130_n 8.52111e-19
cc_20 N_VDD_c_20_p N_VSS_c_130_n 3.48267e-19
cc_21 N_VDD_c_21_p N_VSS_c_134_n 9.21268e-19
cc_22 N_VDD_c_12_p N_VSS_c_134_n 0.00141228f
cc_23 N_VDD_c_4_p N_VSS_c_134_n 0.00225084f
cc_24 N_VDD_c_24_p N_VSS_c_134_n 3.48267e-19
cc_25 N_VDD_XI3.X0_S N_VSS_c_138_n 2.35318e-19
cc_26 N_VDD_c_26_p N_VSS_c_138_n 2.72094e-19
cc_27 N_VDD_c_9_p N_VSS_c_138_n 0.00534617f
cc_28 N_VDD_c_4_p N_VSS_c_138_n 4.25159e-19
cc_29 N_VDD_c_20_p N_VSS_c_138_n 9.58524e-19
cc_30 N_VDD_XI7.X0_S N_VSS_c_143_n 2.15082e-19
cc_31 N_VDD_c_7_p N_VSS_c_143_n 3.16299e-19
cc_32 N_VDD_c_17_p N_VSS_c_145_n 3.66936e-19
cc_33 N_VDD_c_9_p N_VSS_c_145_n 0.00112249f
cc_34 N_VDD_c_19_p N_VSS_c_145_n 3.99794e-19
cc_35 N_VDD_c_20_p N_VSS_c_145_n 8.03027e-19
cc_36 N_VDD_c_21_p N_VSS_c_149_n 3.82294e-19
cc_37 N_VDD_c_12_p N_VSS_c_149_n 0.00112249f
cc_38 N_VDD_c_4_p N_VSS_c_149_n 9.55322e-19
cc_39 N_VDD_c_24_p N_VSS_c_149_n 8.0279e-19
cc_40 N_VDD_c_17_p N_VSS_c_153_n 0.00287902f
cc_41 N_VDD_c_14_p N_VSS_c_153_n 0.0057117f
cc_42 N_VDD_c_42_p N_VSS_c_153_n 0.0010706f
cc_43 N_VDD_c_14_p N_VSS_c_156_n 0.00304013f
cc_44 N_VDD_c_9_p N_VSS_c_157_n 0.00342836f
cc_45 N_VDD_c_45_p N_VSS_c_158_n 0.00107429f
cc_46 N_VDD_c_16_p N_VSS_c_159_n 0.00352516f
cc_47 N_VDD_c_12_p N_VSS_c_159_n 0.0060405f
cc_48 N_VDD_c_48_p N_VSS_c_159_n 0.00101104f
cc_49 N_VDD_c_49_p N_VSS_c_162_n 0.00105833f
cc_50 N_VDD_c_9_p N_VSS_c_163_n 0.00458401f
cc_51 N_VDD_c_7_p N_VSS_c_164_n 0.00135143f
cc_52 N_VDD_c_14_p N_VSS_c_165_n 7.88896e-19
cc_53 N_VDD_c_9_p N_VSS_c_166_n 7.74609e-19
cc_54 N_VDD_c_4_p N_A_XI8.X0_PGD 2.51969e-19
cc_55 N_VDD_c_24_p N_A_c_214_n 0.00237738f
cc_56 N_VDD_XI9.X0_PGD N_A_c_215_n 4.04053e-19
cc_57 N_VDD_XI10.X0_PGD N_A_c_215_n 2.40582e-19
cc_58 N_VDD_c_58_p N_A_c_217_n 9.54306e-19
cc_59 N_VDD_XI10.X0_PGD N_A_c_218_n 2.40582e-19
cc_60 N_VDD_c_60_p N_A_c_219_n 5.838e-19
cc_61 N_VDD_c_14_p N_A_c_220_n 5.24876e-19
cc_62 N_VDD_c_21_p N_A_c_220_n 6.41525e-19
cc_63 N_VDD_c_24_p N_A_c_220_n 4.56568e-19
cc_64 N_VDD_c_4_p N_A_c_223_n 0.00237851f
cc_65 N_VDD_c_60_p N_A_c_223_n 0.00200281f
cc_66 N_VDD_c_60_p N_A_c_225_n 8.17097e-19
cc_67 N_VDD_c_14_p N_A_c_226_n 6.27972e-19
cc_68 N_VDD_c_21_p N_A_c_226_n 4.85469e-19
cc_69 N_VDD_c_24_p N_A_c_226_n 6.1245e-19
cc_70 N_VDD_c_4_p N_A_c_229_n 9.84209e-19
cc_71 N_VDD_c_60_p N_A_c_229_n 2.37583e-19
cc_72 N_VDD_XI1.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_73 N_VDD_c_9_p N_NET1_XI1.X0_D 3.7884e-19
cc_74 N_VDD_c_3_p N_NET1_XI1.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_S N_NET1_c_276_n 3.48267e-19
cc_76 N_VDD_c_9_p N_NET1_c_276_n 4.58491e-19
cc_77 N_VDD_c_3_p N_NET1_c_276_n 5.226e-19
cc_78 N_VDD_c_19_p N_NET1_c_279_n 0.00121121f
cc_79 N_VDD_c_9_p N_NET1_c_280_n 3.78572e-19
cc_80 N_VDD_XI3.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_81 N_VDD_c_12_p N_NET2_XI9.X0_D 3.7884e-19
cc_82 N_VDD_c_4_p N_NET2_XI9.X0_D 3.48267e-19
cc_83 N_VDD_c_60_p N_NET2_c_314_n 8.01015e-19
cc_84 N_VDD_XI3.X0_S N_NET2_c_315_n 3.48267e-19
cc_85 N_VDD_c_12_p N_NET2_c_315_n 4.58491e-19
cc_86 N_VDD_c_4_p N_NET2_c_315_n 8.45449e-19
cc_87 N_VDD_c_12_p N_NET2_c_318_n 3.29894e-19
cc_88 N_VDD_c_4_p N_NET2_c_318_n 8.51778e-19
cc_89 N_VDD_c_60_p N_NET2_c_318_n 0.00334727f
cc_90 N_VDD_c_90_p N_NET2_c_318_n 7.7731e-19
cc_91 N_VDD_c_60_p N_NET2_c_322_n 2.33029e-19
cc_92 N_VDD_c_90_p N_NET2_c_322_n 3.66936e-19
cc_93 N_VDD_c_21_p N_NET2_c_324_n 3.10284e-19
cc_94 N_VDD_c_20_p N_B_XI10.X0_CG 0.00237871f
cc_95 N_VDD_XI10.X0_PGD N_B_XI5.X0_PGD 0.00176522f
cc_96 N_VDD_XI9.X0_PGD N_B_c_363_n 2.40582e-19
cc_97 N_VDD_XI10.X0_PGD N_B_c_363_n 4.04053e-19
cc_98 N_VDD_XI10.X0_PGD N_B_c_365_n 4.05198e-19
cc_99 N_VDD_c_26_p N_B_c_366_n 0.00154836f
cc_100 N_VDD_c_19_p N_B_c_367_n 5.50671e-19
cc_101 N_VDD_c_20_p N_B_c_367_n 8.9014e-19
cc_102 N_VDD_c_19_p N_B_c_369_n 4.73723e-19
cc_103 N_VDD_c_20_p N_B_c_369_n 0.0014909f
cc_104 N_VDD_XI3.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_105 N_VDD_XI7.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_106 N_VDD_c_4_p N_Z_XI8.X0_D 3.48267e-19
cc_107 N_VDD_c_60_p N_Z_XI8.X0_D 3.7884e-19
cc_108 N_VDD_c_7_p N_Z_XI8.X0_D 3.72199e-19
cc_109 N_VDD_XI3.X0_S N_Z_c_403_n 3.48267e-19
cc_110 N_VDD_XI7.X0_S N_Z_c_403_n 3.48267e-19
cc_111 N_VDD_c_4_p N_Z_c_403_n 5.21254e-19
cc_112 N_VDD_c_60_p N_Z_c_403_n 6.55718e-19
cc_113 N_VDD_c_7_p N_Z_c_403_n 8.25922e-19
cc_114 N_VSS_c_149_n N_A_XI3.X0_CG 9.02944e-19
cc_115 N_VSS_XI3.X0_PGD N_A_XI8.X0_PGD 0.00150976f
cc_116 N_VSS_XI1.X0_PGD N_A_c_215_n 2.40582e-19
cc_117 N_VSS_XI3.X0_PGD N_A_c_215_n 3.99472e-19
cc_118 N_VSS_XI3.X0_PGD N_A_c_218_n 4.05198e-19
cc_119 N_VSS_c_172_p N_A_c_219_n 0.00150976f
cc_120 N_VSS_c_134_n N_A_c_223_n 4.12959e-19
cc_121 N_VSS_c_153_n N_A_c_223_n 3.96361e-19
cc_122 N_VSS_c_163_n N_A_c_225_n 2.41875e-19
cc_123 N_VSS_c_145_n N_A_c_226_n 4.65658e-19
cc_124 N_VSS_c_149_n N_A_c_229_n 8.90609e-19
cc_125 N_VSS_c_163_n N_A_c_242_n 3.10545e-19
cc_126 N_VSS_XI10.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_127 N_VSS_c_138_n N_NET1_XI1.X0_D 3.48267e-19
cc_128 N_VSS_XI10.X0_S N_NET1_c_276_n 3.48267e-19
cc_129 N_VSS_c_138_n N_NET1_c_276_n 0.0012813f
cc_130 N_VSS_c_138_n N_NET1_c_279_n 0.00174104f
cc_131 N_VSS_c_163_n N_NET1_c_279_n 5.89244e-19
cc_132 N_VSS_c_185_p N_NET1_c_279_n 0.00121599f
cc_133 N_VSS_c_130_n N_NET1_c_280_n 0.00206231f
cc_134 N_VSS_c_153_n N_NET1_c_280_n 9.32604e-19
cc_135 N_VSS_c_163_n N_NET1_c_280_n 0.0214545f
cc_136 N_VSS_XI9.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_137 N_VSS_c_126_n N_NET2_XI9.X0_D 3.48267e-19
cc_138 N_VSS_XI9.X0_S N_NET2_c_315_n 3.48267e-19
cc_139 N_VSS_c_126_n N_NET2_c_315_n 0.00108327f
cc_140 N_VSS_c_159_n N_NET2_c_315_n 3.31434e-19
cc_141 N_VSS_c_134_n N_NET2_c_318_n 0.00143089f
cc_142 N_VSS_c_156_n N_NET2_c_324_n 3.36104e-19
cc_143 N_VSS_c_159_n N_NET2_c_324_n 6.48614e-19
cc_144 N_VSS_c_145_n N_B_XI1.X0_CG 9.02944e-19
cc_145 N_VSS_XI1.X0_PGD N_B_c_363_n 3.99472e-19
cc_146 N_VSS_XI3.X0_PGD N_B_c_363_n 2.40582e-19
cc_147 N_VSS_XI3.X0_PGD N_B_c_365_n 2.40582e-19
cc_148 N_VSS_c_138_n N_B_c_366_n 2.8419e-19
cc_149 N_VSS_c_149_n N_B_c_367_n 2.07877e-19
cc_150 N_VSS_c_153_n N_B_c_367_n 2.27769e-19
cc_151 N_VSS_c_149_n N_B_c_369_n 7.33679e-19
cc_152 N_VSS_XI10.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_153 N_VSS_XI11.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_154 N_VSS_c_138_n N_Z_XI5.X0_D 3.48267e-19
cc_155 N_VSS_c_143_n N_Z_XI5.X0_D 3.48267e-19
cc_156 N_VSS_XI10.X0_S N_Z_c_403_n 3.48267e-19
cc_157 N_VSS_XI11.X0_S N_Z_c_403_n 3.48267e-19
cc_158 N_VSS_c_138_n N_Z_c_403_n 8.61925e-19
cc_159 N_VSS_c_143_n N_Z_c_403_n 5.69026e-19
cc_160 N_A_XI11.X0_CG N_NET1_XI11.X0_PGD 4.5346e-19
cc_161 N_A_c_244_p N_NET1_XI11.X0_PGD 0.00151381f
cc_162 N_A_c_244_p N_NET1_c_293_n 0.00157635f
cc_163 N_A_c_225_n N_NET1_c_279_n 0.00310276f
cc_164 N_A_c_242_n N_NET1_c_279_n 0.00205512f
cc_165 N_A_XI11.X0_CG N_NET1_c_296_n 0.00234108f
cc_166 N_A_c_249_p N_NET1_c_296_n 0.00101616f
cc_167 N_A_c_244_p N_NET1_c_296_n 0.00161406f
cc_168 N_A_XI8.X0_PGD N_NET2_XI7.X0_PGD 0.00160287f
cc_169 N_A_c_218_n N_NET2_XI7.X0_PGD 3.14428e-19
cc_170 N_A_c_244_p N_NET2_XI7.X0_PGD 5.68075e-19
cc_171 N_A_XI8.X0_PGD N_NET2_c_336_n 4.60549e-19
cc_172 N_A_c_219_n N_NET2_c_314_n 0.00160287f
cc_173 N_A_c_223_n N_NET2_c_315_n 7.37727e-19
cc_174 N_A_c_223_n N_NET2_c_318_n 0.00205074f
cc_175 N_A_c_225_n N_NET2_c_318_n 0.0018485f
cc_176 N_A_c_229_n N_NET2_c_318_n 3.44698e-19
cc_177 N_A_c_223_n N_NET2_c_322_n 3.44698e-19
cc_178 N_A_c_229_n N_NET2_c_322_n 9.07485e-19
cc_179 N_A_c_244_p N_NET2_c_322_n 3.98239e-19
cc_180 N_A_c_218_n N_B_XI8.X0_CG 0.003858f
cc_181 N_A_c_229_n N_B_XI8.X0_CG 0.00111269f
cc_182 N_A_c_215_n N_B_c_363_n 0.00575421f
cc_183 N_A_c_226_n N_B_c_382_n 4.09767e-19
cc_184 N_A_c_218_n N_B_c_365_n 0.00308843f
cc_185 N_A_c_218_n N_B_c_384_n 0.00362155f
cc_186 N_A_c_215_n N_B_c_369_n 6.77269e-19
cc_187 N_A_c_223_n N_Z_c_403_n 0.00321233f
cc_188 N_A_c_225_n N_Z_c_403_n 0.0025035f
cc_189 N_A_c_244_p N_Z_c_403_n 8.50872e-19
cc_190 N_NET1_c_276_n N_NET2_XI9.X0_D 2.15082e-19
cc_191 N_NET1_XI11.X0_PGD N_NET2_XI5.X0_CG 2.62058e-19
cc_192 N_NET1_c_293_n N_NET2_XI7.X0_PGD 0.00832016f
cc_193 N_NET1_XI11.X0_PGD N_NET2_c_336_n 0.00416722f
cc_194 N_NET1_XI1.X0_D N_NET2_c_315_n 2.15082e-19
cc_195 N_NET1_c_279_n N_NET2_c_318_n 0.00142494f
cc_196 N_NET1_XI7.X0_CG N_NET2_c_322_n 0.00102831f
cc_197 N_NET1_XI11.X0_PGD N_B_XI5.X0_PGD 0.00188492f
cc_198 N_NET1_XI7.X0_CG N_B_XI8.X0_CG 2.60667e-19
cc_199 N_NET1_c_293_n N_B_c_388_n 2.60667e-19
cc_200 N_NET1_c_309_p N_B_c_366_n 0.00165894f
cc_201 N_NET1_c_279_n N_Z_c_403_n 3.02205e-19
cc_202 N_NET2_XI5.X0_CG N_B_XI5.X0_PGD 0.0019183f
cc_203 N_NET2_c_336_n N_B_XI5.X0_PGD 0.00161994f
cc_204 N_NET2_XI7.X0_PGD N_B_c_392_n 3.1641e-19
cc_205 N_NET2_XI7.X0_PGD N_B_c_388_n 0.00313953f
cc_206 N_NET2_c_356_p N_B_c_388_n 0.00172424f
cc_207 N_NET2_c_356_p N_B_c_395_n 0.0019183f
cc_208 N_NET2_XI7.X0_PGD N_Z_c_403_n 0.00115814f
cc_209 N_NET2_c_336_n N_Z_c_403_n 5.21666e-19
cc_210 N_NET2_c_318_n N_Z_c_403_n 2.80086e-19
cc_211 N_B_c_388_n N_Z_c_403_n 8.84927e-19
cc_212 N_B_c_367_n N_Z_c_403_n 3.17615e-19
*
.ends
*
*
.subckt XNOR2_HPNW1 A B Y VDD VSS
xgate (VDD VSS A B Y) G4_XNOR2_N1
.ends
*
* File: G5_XNOR3_N1.pex.netlist
* Created: Fri Mar 25 15:42:00 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XNOR3_N1_VDD 2 5 9 12 14 17 34 35 44 45 54 55 77 79 80 81 84 86 90
+ 93 96 98 102 104 108 112 114 116 118 119 125 134 139 Vss
c122 139 Vss 0.00481852f
c123 134 Vss 0.00580927f
c124 125 Vss 0.00558883f
c125 119 Vss 2.39889e-19
c126 118 Vss 4.91159e-19
c127 117 Vss 4.14624e-19
c128 114 Vss 3.56526e-19
c129 112 Vss 0.00104518f
c130 108 Vss 3.94646e-19
c131 104 Vss 0.00602085f
c132 102 Vss 0.00109141f
c133 98 Vss 0.00553212f
c134 96 Vss 0.0016276f
c135 93 Vss 0.00243759f
c136 90 Vss 0.00352468f
c137 86 Vss 0.00659816f
c138 84 Vss 0.0015095f
c139 81 Vss 8.67152e-19
c140 80 Vss 0.00945954f
c141 79 Vss 0.00914208f
c142 77 Vss 0.00176824f
c143 57 Vss 5.45153e-20
c144 55 Vss 0.0336444f
c145 54 Vss 0.0988545f
c146 45 Vss 0.0346156f
c147 44 Vss 0.1003f
c148 35 Vss 0.0346129f
c149 34 Vss 0.0990563f
c150 17 Vss 0.165098f
c151 14 Vss 0.00210084f
c152 12 Vss 0.00231756f
c153 9 Vss 0.16518f
c154 5 Vss 0.165156f
c155 2 Vss 0.00208065f
r156 110 112 4.83471
r157 108 139 1.16709
r158 106 108 2.16729
r159 105 119 0.494161
r160 104 110 0.652036
r161 104 105 7.46046
r162 102 134 1.16709
r163 100 119 0.128424
r164 100 102 2.16729
r165 99 118 0.494161
r166 98 106 0.652036
r167 98 99 10.3363
r168 94 117 0.0828784
r169 94 96 2.00578
r170 93 118 0.128424
r171 92 117 0.551426
r172 92 93 4.16786
r173 90 125 1.16709
r174 88 117 0.551426
r175 88 90 5.835
r176 87 116 0.326018
r177 86 118 0.494161
r178 86 87 10.1279
r179 82 114 0.0828784
r180 82 84 1.82344
r181 80 119 0.494161
r182 80 81 15.8795
r183 79 116 0.326018
r184 78 114 0.551426
r185 78 79 13.3371
r186 77 114 0.551426
r187 76 81 0.652036
r188 76 77 4.16786
r189 57 139 0.238214
r190 55 57 1.45875
r191 54 58 0.652036
r192 54 57 1.45875
r193 51 55 0.652036
r194 47 134 0.238214
r195 45 47 1.45875
r196 44 48 0.652036
r197 44 47 1.45875
r198 41 45 0.652036
r199 37 125 0.238214
r200 35 37 1.45875
r201 34 38 0.652036
r202 34 37 1.45875
r203 31 35 0.652036
r204 17 58 2.5674
r205 17 51 2.5674
r206 14 112 1.16709
r207 12 96 1.16709
r208 9 48 2.5674
r209 9 41 2.5674
r210 5 38 2.5674
r211 5 31 2.5674
r212 2 84 1.16709
.ends

.subckt PM_G5_XNOR3_N1_C 2 4 6 8 17 20 23 40 43 47 52 57 62 85 87 93 98 Vss
c60 98 Vss 8.02961e-19
c61 93 Vss 6.27504e-19
c62 87 Vss 0.0049214f
c63 85 Vss 0.00877979f
c64 62 Vss 0.00258187f
c65 57 Vss 0.00458232f
c66 52 Vss 0.00201471f
c67 47 Vss 4.03464e-19
c68 43 Vss 3.73849e-19
c69 40 Vss 5.60764e-19
c70 23 Vss 1.05295e-19
c71 20 Vss 0.220565f
c72 17 Vss 0.0715834f
c73 15 Vss 0.0247918f
c74 8 Vss 0.00236553f
c75 4 Vss 0.0826049f
r76 88 98 0.0685365
r77 87 89 0.652036
r78 87 88 10.3363
r79 86 93 0.0685365
r80 85 98 0.0685365
r81 85 86 24.7154
r82 52 89 2.16729
r83 47 62 1.16709
r84 47 98 2.12561
r85 43 57 1.16709
r86 43 93 0.5835
r87 40 43 0.0416786
r88 23 57 0.0476429
r89 21 23 0.326018
r90 21 23 0.1167
r91 20 24 0.652036
r92 20 23 6.7686
r93 17 57 0.357321
r94 15 23 0.326018
r95 15 17 0.40845
r96 8 52 1.16709
r97 6 62 0.75
r98 4 24 2.5674
r99 2 17 2.15895
.ends

.subckt PM_G5_XNOR3_N1_VSS 3 6 11 15 18 34 37 44 45 47 54 55 73 78 83 88 93 96
+ 99 108 113 122 124 125 126 131 132 137 145 153 154 155 Vss
c131 155 Vss 3.75522e-19
c132 154 Vss 3.87529e-19
c133 153 Vss 4.4306e-19
c134 137 Vss 0.00333207f
c135 132 Vss 8.38361e-19
c136 131 Vss 0.00578307f
c137 126 Vss 8.35423e-19
c138 125 Vss 0.00509728f
c139 124 Vss 0.0036146f
c140 122 Vss 0.00254978f
c141 113 Vss 0.00381203f
c142 108 Vss 0.0040091f
c143 99 Vss 0.00484046f
c144 96 Vss 0.00348301f
c145 93 Vss 0.00279856f
c146 88 Vss 7.12901e-19
c147 83 Vss 0.00141291f
c148 78 Vss 0.0025656f
c149 73 Vss 0.00249897f
c150 55 Vss 0.0338093f
c151 54 Vss 0.0988897f
c152 47 Vss 7.60188e-20
c153 45 Vss 0.0331638f
c154 44 Vss 0.0974849f
c155 37 Vss 7.50699e-20
c156 35 Vss 0.0349827f
c157 34 Vss 0.1003f
c158 18 Vss 0.00263959f
c159 15 Vss 0.164604f
c160 11 Vss 0.166952f
c161 6 Vss 0.00172036f
c162 3 Vss 0.167004f
r163 143 155 0.494161
r164 143 145 6.71025
r165 139 155 0.128424
r166 138 154 0.494161
r167 137 149 0.652036
r168 137 138 7.46046
r169 133 154 0.128424
r170 131 155 0.494161
r171 131 132 15.8795
r172 127 153 0.0828784
r173 125 154 0.494161
r174 125 126 13.0037
r175 124 132 0.652036
r176 123 153 0.551426
r177 123 124 10.6697
r178 122 153 0.551426
r179 121 126 0.652036
r180 121 122 6.83529
r181 96 145 1.33371
r182 93 96 5.41821
r183 88 113 1.16709
r184 88 149 2.16729
r185 83 108 1.16709
r186 83 139 2.16729
r187 78 133 4.83471
r188 73 99 1.16709
r189 73 127 4.33978
r190 57 113 0.238214
r191 55 57 1.45875
r192 54 58 0.652036
r193 54 57 1.45875
r194 51 55 0.652036
r195 47 108 0.238214
r196 45 47 1.45875
r197 44 48 0.652036
r198 44 47 1.45875
r199 41 45 0.652036
r200 37 99 0.238214
r201 35 37 1.45875
r202 34 38 0.652036
r203 34 37 1.45875
r204 31 35 0.652036
r205 18 93 1.16709
r206 15 58 2.5674
r207 15 51 2.5674
r208 11 48 2.5674
r209 11 41 2.5674
r210 6 78 1.16709
r211 3 38 2.5674
r212 3 31 2.5674
.ends

.subckt PM_G5_XNOR3_N1_CI 2 6 8 34 39 44 79 80 85 91 Vss
c47 91 Vss 2.52123e-19
c48 85 Vss 0.00547442f
c49 80 Vss 3.74154e-19
c50 79 Vss 0.0039666f
c51 44 Vss 0.00209085f
c52 39 Vss 0.00132824f
c53 34 Vss 0.00535743f
c54 8 Vss 0.00276539f
c55 6 Vss 0.00213002f
c56 2 Vss 0.00154503f
r57 86 91 0.494161
r58 85 87 0.652036
r59 85 86 10.3363
r60 81 91 0.128424
r61 79 91 0.494161
r62 79 80 21.8396
r63 75 80 0.652036
r64 44 87 2.16729
r65 39 81 2.16729
r66 34 75 11.3366
r67 8 44 1.16709
r68 6 39 1.16709
r69 2 34 1.16709
.ends

.subckt PM_G5_XNOR3_N1_A 2 4 7 11 21 24 45 49 51 54 56 57 58 62 63 69 74 Vss
c79 74 Vss 0.00491901f
c80 69 Vss 0.00491594f
c81 63 Vss 8.26639e-19
c82 62 Vss 4.20301e-19
c83 58 Vss 0.0011362f
c84 57 Vss 0.00976615f
c85 56 Vss 0.00370619f
c86 51 Vss 0.00520175f
c87 49 Vss 0.135015f
c88 45 Vss 0.126353f
c89 24 Vss 0.2139f
c90 21 Vss 0.0724995f
c91 19 Vss 0.0247918f
c92 7 Vss 1.00425f
c93 4 Vss 0.0850321f
r94 74 77 0.1
r95 66 77 1.16709
r96 63 66 0.833571
r97 60 69 1.16709
r98 60 62 0.513084
r99 57 63 0.0685365
r100 57 58 10.4613
r101 55 58 0.652036
r102 55 56 8.66914
r103 54 62 0.791893
r104 51 56 0.652036
r105 51 54 9.41936
r106 47 49 4.53833
r107 44 74 0.262036
r108 44 45 2.26917
r109 41 44 2.26917
r110 36 49 0.00605528
r111 35 45 0.00605528
r112 32 47 0.00605528
r113 31 41 0.00605528
r114 27 69 0.0952857
r115 25 27 0.326018
r116 25 27 0.1167
r117 24 28 0.652036
r118 24 27 6.7686
r119 21 27 0.3335
r120 19 27 0.326018
r121 19 21 0.2334
r122 11 36 2.5674
r123 11 32 2.5674
r124 7 11 12.837
r125 7 35 2.5674
r126 7 11 12.837
r127 7 31 2.5674
r128 4 28 2.5674
r129 2 21 2.334
.ends

.subckt PM_G5_XNOR3_N1_BI 2 6 8 16 23 32 37 42 51 56 64 65 71 78 83 84 Vss
c70 84 Vss 1.10364e-19
c71 83 Vss 0.00214683f
c72 78 Vss 8.34553e-19
c73 71 Vss 5.02505e-19
c74 65 Vss 4.43116e-19
c75 64 Vss 0.00191151f
c76 56 Vss 0.00250766f
c77 51 Vss 0.00202351f
c78 42 Vss 0.00122467f
c79 37 Vss 4.09629e-19
c80 32 Vss 0.00157267f
c81 23 Vss 7.03109e-20
c82 16 Vss 0.0573997f
c83 8 Vss 0.0573997f
c84 2 Vss 0.00150258f
r85 82 84 0.65228
r86 82 83 3.46076
r87 78 83 0.65228
r88 74 78 2.1006
r89 71 74 2.08393
r90 64 71 0.0685365
r91 64 65 13.2121
r92 60 65 0.652036
r93 42 56 1.16709
r94 42 84 2.1395
r95 37 51 1.16709
r96 37 74 0.0416786
r97 32 60 4.29289
r98 23 56 0.50025
r99 16 51 0.50025
r100 8 23 1.80885
r101 6 16 1.80885
r102 2 32 1.16709
.ends

.subckt PM_G5_XNOR3_N1_AI 2 7 11 31 36 37 46 51 60 69 Vss
c47 69 Vss 2.92061e-19
c48 60 Vss 0.0055297f
c49 51 Vss 0.00389112f
c50 46 Vss 9.98085e-19
c51 37 Vss 0.127837f
c52 36 Vss 5.86204e-20
c53 31 Vss 0.128631f
c54 7 Vss 0.994815f
c55 2 Vss 0.00150258f
r56 65 69 0.652036
r57 60 63 0.1
r58 51 63 1.16709
r59 51 69 13.7539
r60 46 65 2.16729
r61 36 60 0.262036
r62 36 37 2.334
r63 33 36 2.20433
r64 29 31 4.53833
r65 26 37 0.00605528
r66 25 31 0.00605528
r67 22 33 0.00605528
r68 21 29 0.00605528
r69 11 26 2.5674
r70 11 22 2.5674
r71 7 11 12.837
r72 7 25 2.5674
r73 7 11 12.837
r74 7 21 2.5674
r75 2 46 1.16709
.ends

.subckt PM_G5_XNOR3_N1_B 2 4 6 8 16 17 24 28 31 42 45 50 55 60 65 69 76 77 Vss
c63 77 Vss 1.47395e-19
c64 76 Vss 6.32207e-19
c65 69 Vss 0.0035022f
c66 65 Vss 0.00265398f
c67 60 Vss 0.00253939f
c68 55 Vss 0.00274111f
c69 50 Vss 0.00171367f
c70 45 Vss 5.45343e-20
c71 42 Vss 5.46775e-19
c72 31 Vss 0.0573997f
c73 24 Vss 1.2014e-19
c74 20 Vss 0.0247918f
c75 17 Vss 0.0338376f
c76 16 Vss 0.183114f
c77 6 Vss 0.0573997f
c78 4 Vss 0.0714101f
c79 2 Vss 0.0826049f
r80 76 77 0.65228
r81 75 76 3.46076
r82 69 75 0.65228
r83 50 65 1.16709
r84 50 77 2.1395
r85 45 60 1.16709
r86 45 69 2.1006
r87 38 55 1.16709
r88 38 45 10.7364
r89 38 42 0.0364688
r90 36 55 0.0476429
r91 31 65 0.50025
r92 28 60 0.50025
r93 24 55 0.357321
r94 20 36 0.326018
r95 20 24 0.40845
r96 17 36 6.7686
r97 16 36 0.326018
r98 16 36 0.1167
r99 13 17 0.652036
r100 8 31 1.80885
r101 6 28 1.80885
r102 4 24 2.15895
r103 2 13 2.5674
.ends

.subckt PM_G5_XNOR3_N1_Z 2 4 30 33 Vss
c31 30 Vss 0.00315811f
c32 4 Vss 0.00153036f
c33 2 Vss 0.00166246f
r34 33 35 4.20954
r35 30 33 4.95975
r36 4 35 1.16709
r37 2 30 1.16709
.ends

.subckt G5_XNOR3_N1  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI10.X0 N_CI_XI10.X0_D N_VSS_XI10.X0_PGD N_C_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW1
XI9.X0 N_CI_XI10.X0_D N_VDD_XI9.X0_PGD N_C_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW1
XI5.X0 N_BI_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW1
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW1
XI6.X0 N_BI_XI5.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW1
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW1
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_B_XI2.X0_CG N_AI_XI2.X0_PGD N_C_XI2.X0_S
+ TIGFET_HPNW1
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_BI_XI4.X0_CG N_AI_XI4.X0_PGD N_CI_XI4.X0_S
+ TIGFET_HPNW1
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_BI_XI3.X0_CG N_A_XI3.X0_PGD N_C_XI3.X0_S
+ TIGFET_HPNW1
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_B_XI1.X0_CG N_A_XI1.X0_PGD N_CI_XI1.X0_S
+ TIGFET_HPNW1
*
x_PM_G5_XNOR3_N1_VDD N_VDD_XI10.X0_S N_VDD_XI9.X0_PGD N_VDD_XI5.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI6.X0_S N_VDD_XI7.X0_PGD N_VDD_c_120_p N_VDD_c_18_p
+ N_VDD_c_23_p N_VDD_c_4_p N_VDD_c_110_p N_VDD_c_19_p N_VDD_c_6_p N_VDD_c_25_p
+ N_VDD_c_5_p N_VDD_c_64_p N_VDD_c_27_p N_VDD_c_28_p N_VDD_c_29_p N_VDD_c_35_p
+ N_VDD_c_32_p N_VDD_c_20_p N_VDD_c_11_p N_VDD_c_24_p N_VDD_c_37_p N_VDD_c_12_p
+ N_VDD_c_60_p VDD N_VDD_c_68_p N_VDD_c_72_p N_VDD_c_2_p N_VDD_c_42_p
+ N_VDD_c_38_p Vss PM_G5_XNOR3_N1_VDD
x_PM_G5_XNOR3_N1_C N_C_XI10.X0_CG N_C_XI9.X0_CG N_C_XI2.X0_S N_C_XI3.X0_S
+ N_C_c_143_p N_C_c_125_n N_C_c_136_p C N_C_c_138_p N_C_c_158_p N_C_c_178_p
+ N_C_c_130_n N_C_c_132_n N_C_c_133_n N_C_c_156_p N_C_c_139_p N_C_c_161_p Vss
+ PM_G5_XNOR3_N1_C
x_PM_G5_XNOR3_N1_VSS N_VSS_XI10.X0_PGD N_VSS_XI9.X0_S N_VSS_XI8.X0_PGD
+ N_VSS_XI6.X0_PGD N_VSS_XI7.X0_S N_VSS_c_188_n N_VSS_c_247_n N_VSS_c_189_n
+ N_VSS_c_191_n N_VSS_c_287_p N_VSS_c_192_n N_VSS_c_193_n N_VSS_c_195_n
+ N_VSS_c_201_n N_VSS_c_205_n N_VSS_c_209_n N_VSS_c_213_n N_VSS_c_216_n
+ N_VSS_c_217_n N_VSS_c_220_n N_VSS_c_224_n N_VSS_c_228_n N_VSS_c_231_n
+ N_VSS_c_233_n N_VSS_c_234_n N_VSS_c_235_n N_VSS_c_239_n N_VSS_c_240_n VSS
+ N_VSS_c_243_n N_VSS_c_244_n N_VSS_c_245_n Vss PM_G5_XNOR3_N1_VSS
x_PM_G5_XNOR3_N1_CI N_CI_XI10.X0_D N_CI_XI4.X0_S N_CI_XI1.X0_S N_CI_c_316_n
+ N_CI_c_334_n N_CI_c_356_p N_CI_c_320_n N_CI_c_338_n N_CI_c_324_n N_CI_c_349_p
+ Vss PM_G5_XNOR3_N1_CI
x_PM_G5_XNOR3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI3.X0_PGD N_A_XI1.X0_PGD
+ N_A_c_387_n N_A_c_362_n N_A_c_415_p N_A_c_417_p N_A_c_363_n A N_A_c_370_n
+ N_A_c_381_n N_A_c_371_n N_A_c_372_n N_A_c_386_n N_A_c_374_n N_A_c_399_p Vss
+ PM_G5_XNOR3_N1_A
x_PM_G5_XNOR3_N1_BI N_BI_XI5.X0_D N_BI_XI4.X0_CG N_BI_XI3.X0_CG N_BI_c_478_p
+ N_BI_c_465_n N_BI_c_443_n N_BI_c_468_n N_BI_c_459_n N_BI_c_471_n N_BI_c_472_n
+ N_BI_c_447_n N_BI_c_457_n N_BI_c_477_n N_BI_c_450_n N_BI_c_503_p N_BI_c_451_n
+ Vss PM_G5_XNOR3_N1_BI
x_PM_G5_XNOR3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_523_n
+ N_AI_c_546_n N_AI_c_513_n N_AI_c_514_n N_AI_c_517_n N_AI_c_528_n N_AI_c_518_n
+ Vss PM_G5_XNOR3_N1_AI
x_PM_G5_XNOR3_N1_B N_B_XI5.X0_CG N_B_XI6.X0_CG N_B_XI2.X0_CG N_B_XI1.X0_CG
+ N_B_c_559_n N_B_c_561_n N_B_c_571_n N_B_c_580_n N_B_c_581_n B N_B_c_584_n
+ N_B_c_575_n N_B_c_562_n N_B_c_589_n N_B_c_590_n N_B_c_563_n N_B_c_607_n
+ N_B_c_576_n Vss PM_G5_XNOR3_N1_B
x_PM_G5_XNOR3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_624_n Z Vss PM_G5_XNOR3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_C_XI9.X0_CG 9.58934e-19
cc_2 N_VDD_c_2_p N_C_XI9.X0_CG 8.03148e-19
cc_3 N_VDD_XI9.X0_PGD N_C_c_125_n 4.16623e-19
cc_4 N_VDD_c_4_p N_C_c_125_n 9.58934e-19
cc_5 N_VDD_c_5_p N_C_c_125_n 0.00125128f
cc_6 N_VDD_c_6_p C 3.00172e-19
cc_7 N_VDD_c_5_p C 0.00118142f
cc_8 N_VDD_c_6_p N_C_c_130_n 4.71537e-19
cc_9 N_VDD_c_5_p N_C_c_130_n 2.74773e-19
cc_10 N_VDD_XI6.X0_S N_C_c_132_n 3.43419e-19
cc_11 N_VDD_c_11_p N_C_c_133_n 5.30636e-19
cc_12 N_VDD_c_12_p N_C_c_133_n 7.99481e-19
cc_13 N_VDD_XI9.X0_PGD N_VSS_XI10.X0_PGD 0.00173038f
cc_14 N_VDD_XI5.X0_PGD N_VSS_XI8.X0_PGD 2.27468e-19
cc_15 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172039f
cc_16 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017188f
cc_17 N_VDD_XI7.X0_PGD N_VSS_XI6.X0_PGD 2.1536e-19
cc_18 N_VDD_c_18_p N_VSS_c_188_n 0.00173038f
cc_19 N_VDD_c_19_p N_VSS_c_189_n 0.00172039f
cc_20 N_VDD_c_20_p N_VSS_c_189_n 2.46461e-19
cc_21 N_VDD_c_20_p N_VSS_c_191_n 3.60588e-19
cc_22 N_VDD_c_12_p N_VSS_c_192_n 2.35445e-19
cc_23 N_VDD_c_23_p N_VSS_c_193_n 0.0017188f
cc_24 N_VDD_c_24_p N_VSS_c_193_n 2.74208e-19
cc_25 N_VDD_c_25_p N_VSS_c_195_n 4.32468e-19
cc_26 N_VDD_c_5_p N_VSS_c_195_n 4.60511e-19
cc_27 N_VDD_c_27_p N_VSS_c_195_n 0.00130521f
cc_28 N_VDD_c_28_p N_VSS_c_195_n 4.50568e-19
cc_29 N_VDD_c_29_p N_VSS_c_195_n 3.98949e-19
cc_30 N_VDD_c_2_p N_VSS_c_195_n 3.48267e-19
cc_31 N_VDD_c_5_p N_VSS_c_201_n 5.01863e-19
cc_32 N_VDD_c_32_p N_VSS_c_201_n 2.14355e-19
cc_33 N_VDD_c_11_p N_VSS_c_201_n 7.9087e-19
cc_34 N_VDD_c_12_p N_VSS_c_201_n 3.30117e-19
cc_35 N_VDD_c_35_p N_VSS_c_205_n 6.99368e-19
cc_36 N_VDD_c_20_p N_VSS_c_205_n 0.00161703f
cc_37 N_VDD_c_37_p N_VSS_c_205_n 8.32098e-19
cc_38 N_VDD_c_38_p N_VSS_c_205_n 3.48267e-19
cc_39 N_VDD_c_11_p N_VSS_c_209_n 6.79271e-19
cc_40 N_VDD_c_24_p N_VSS_c_209_n 0.00161703f
cc_41 N_VDD_c_12_p N_VSS_c_209_n 0.00241473f
cc_42 N_VDD_c_42_p N_VSS_c_209_n 3.48267e-19
cc_43 N_VDD_XI7.X0_PGD N_VSS_c_213_n 3.41313e-19
cc_44 N_VDD_c_37_p N_VSS_c_213_n 0.00506009f
cc_45 N_VDD_c_38_p N_VSS_c_213_n 9.58524e-19
cc_46 N_VDD_c_20_p N_VSS_c_216_n 0.00415364f
cc_47 N_VDD_c_25_p N_VSS_c_217_n 4.41003e-19
cc_48 N_VDD_c_29_p N_VSS_c_217_n 3.89161e-19
cc_49 N_VDD_c_2_p N_VSS_c_217_n 7.99831e-19
cc_50 N_VDD_c_35_p N_VSS_c_220_n 3.48267e-19
cc_51 N_VDD_c_20_p N_VSS_c_220_n 2.03837e-19
cc_52 N_VDD_c_37_p N_VSS_c_220_n 3.99794e-19
cc_53 N_VDD_c_38_p N_VSS_c_220_n 8.03027e-19
cc_54 N_VDD_c_11_p N_VSS_c_224_n 3.82294e-19
cc_55 N_VDD_c_24_p N_VSS_c_224_n 2.03837e-19
cc_56 N_VDD_c_12_p N_VSS_c_224_n 9.55109e-19
cc_57 N_VDD_c_42_p N_VSS_c_224_n 8.01441e-19
cc_58 N_VDD_c_6_p N_VSS_c_228_n 0.00301593f
cc_59 N_VDD_c_25_p N_VSS_c_228_n 7.60301e-19
cc_60 N_VDD_c_60_p N_VSS_c_228_n 0.0010705f
cc_61 N_VDD_c_25_p N_VSS_c_231_n 0.00803422f
cc_62 N_VDD_c_29_p N_VSS_c_231_n 8.94414e-19
cc_63 N_VDD_c_5_p N_VSS_c_233_n 0.00969041f
cc_64 N_VDD_c_64_p N_VSS_c_234_n 0.00107143f
cc_65 N_VDD_c_28_p N_VSS_c_235_n 0.00807788f
cc_66 N_VDD_c_32_p N_VSS_c_235_n 7.22996e-19
cc_67 N_VDD_c_20_p N_VSS_c_235_n 0.00374557f
cc_68 N_VDD_c_68_p N_VSS_c_235_n 0.00137227f
cc_69 N_VDD_c_25_p N_VSS_c_239_n 0.00107355f
cc_70 N_VDD_c_5_p N_VSS_c_240_n 0.00142851f
cc_71 N_VDD_c_24_p N_VSS_c_240_n 0.00577339f
cc_72 N_VDD_c_72_p N_VSS_c_240_n 0.00106333f
cc_73 N_VDD_c_25_p N_VSS_c_243_n 0.00112682f
cc_74 N_VDD_c_5_p N_VSS_c_244_n 0.00104966f
cc_75 N_VDD_c_20_p N_VSS_c_245_n 7.74609e-19
cc_76 N_VDD_XI10.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_77 N_VDD_c_27_p N_CI_XI10.X0_D 3.72199e-19
cc_78 N_VDD_XI10.X0_S N_CI_c_316_n 3.48267e-19
cc_79 N_VDD_c_5_p N_CI_c_316_n 5.01863e-19
cc_80 N_VDD_c_27_p N_CI_c_316_n 5.226e-19
cc_81 N_VDD_c_29_p N_CI_c_316_n 0.00213742f
cc_82 N_VDD_c_35_p N_CI_c_320_n 7.47076e-19
cc_83 N_VDD_c_32_p N_CI_c_320_n 4.06004e-19
cc_84 N_VDD_c_38_p N_A_XI7.X0_CG 9.92565e-19
cc_85 N_VDD_XI7.X0_PGD N_A_c_362_n 3.90792e-19
cc_86 N_VDD_XI6.X0_S N_A_c_363_n 2.96819e-19
cc_87 N_VDD_XI7.X0_PGD N_A_c_363_n 5.17967e-19
cc_88 N_VDD_c_20_p N_A_c_363_n 4.32724e-19
cc_89 N_VDD_c_24_p N_A_c_363_n 4.10602e-19
cc_90 N_VDD_c_37_p N_A_c_363_n 4.1682e-19
cc_91 N_VDD_c_12_p N_A_c_363_n 3.91173e-19
cc_92 N_VDD_c_38_p N_A_c_363_n 5.53168e-19
cc_93 N_VDD_XI6.X0_S N_A_c_370_n 9.18655e-19
cc_94 N_VDD_c_12_p N_A_c_371_n 0.00608947f
cc_95 N_VDD_c_29_p N_A_c_372_n 8.16868e-19
cc_96 N_VDD_c_11_p N_A_c_372_n 2.36389e-19
cc_97 N_VDD_c_29_p N_A_c_374_n 6.33536e-19
cc_98 N_VDD_c_42_p N_A_c_374_n 5.39283e-19
cc_99 N_VDD_XI6.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_100 N_VDD_c_24_p N_BI_XI5.X0_D 3.7884e-19
cc_101 N_VDD_c_12_p N_BI_XI5.X0_D 3.48267e-19
cc_102 N_VDD_XI6.X0_S N_BI_c_443_n 3.48267e-19
cc_103 N_VDD_c_29_p N_BI_c_443_n 8.52765e-19
cc_104 N_VDD_c_24_p N_BI_c_443_n 4.58491e-19
cc_105 N_VDD_c_12_p N_BI_c_443_n 7.03408e-19
cc_106 N_VDD_c_24_p N_BI_c_447_n 2.4324e-19
cc_107 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_108 N_VDD_c_32_p N_AI_XI8.X0_D 3.73302e-19
cc_109 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.86706e-19
cc_110 N_VDD_c_110_p N_AI_c_513_n 2.86706e-19
cc_111 N_VDD_XI8.X0_S N_AI_c_514_n 3.48267e-19
cc_112 N_VDD_c_32_p N_AI_c_514_n 5.23123e-19
cc_113 N_VDD_c_20_p N_AI_c_514_n 5.01863e-19
cc_114 N_VDD_c_37_p N_AI_c_517_n 0.00111556f
cc_115 N_VDD_c_20_p N_AI_c_518_n 2.2965e-19
cc_116 N_VDD_XI9.X0_PGD N_B_XI5.X0_CG 9.5906e-19
cc_117 N_VDD_c_42_p N_B_XI5.X0_CG 9.74645e-19
cc_118 N_VDD_XI5.X0_PGD N_B_c_559_n 3.9688e-19
cc_119 N_VDD_XI7.X0_PGD N_B_c_559_n 2.07132e-19
cc_120 N_VDD_c_120_p N_B_c_561_n 9.5906e-19
cc_121 N_VDD_c_38_p N_B_c_562_n 2.92921e-19
cc_122 N_VDD_c_12_p N_B_c_563_n 5.34599e-19
cc_123 N_C_c_125_n N_VSS_XI10.X0_PGD 4.16623e-19
cc_124 N_C_c_136_p N_VSS_c_247_n 9.33417e-19
cc_125 C N_VSS_c_195_n 6.06998e-19
cc_126 N_C_c_138_p N_VSS_c_195_n 4.82229e-19
cc_127 N_C_c_139_p N_VSS_c_195_n 2.78014e-19
cc_128 N_C_c_138_p N_VSS_c_201_n 2.30642e-19
cc_129 N_C_c_133_n N_VSS_c_201_n 0.00197293f
cc_130 N_C_c_133_n N_VSS_c_209_n 0.00165406f
cc_131 N_C_c_143_p N_VSS_c_217_n 0.0041205f
cc_132 N_C_c_136_p N_VSS_c_217_n 7.00195e-19
cc_133 C N_VSS_c_217_n 4.56568e-19
cc_134 N_C_c_130_n N_VSS_c_217_n 6.1245e-19
cc_135 C N_VSS_c_228_n 2.17246e-19
cc_136 N_C_c_138_p N_VSS_c_228_n 4.01014e-19
cc_137 N_C_c_139_p N_VSS_c_228_n 4.34874e-19
cc_138 C N_VSS_c_233_n 2.70819e-19
cc_139 N_C_c_138_p N_VSS_c_233_n 9.65301e-19
cc_140 N_C_c_139_p N_VSS_c_233_n 0.00282977f
cc_141 N_C_c_133_n N_VSS_c_240_n 0.00175198f
cc_142 N_C_c_133_n N_CI_c_316_n 0.00136327f
cc_143 N_C_c_133_n N_CI_c_320_n 0.00242327f
cc_144 N_C_c_156_p N_CI_c_324_n 4.1018e-19
cc_145 N_C_c_133_n N_A_c_363_n 2.5075e-19
cc_146 N_C_c_158_p N_A_c_370_n 0.00148519f
cc_147 N_C_c_132_n N_A_c_370_n 8.20481e-19
cc_148 N_C_c_133_n N_A_c_370_n 2.96346e-19
cc_149 N_C_c_161_p N_A_c_370_n 2.4205e-19
cc_150 N_C_c_158_p N_A_c_381_n 0.00189731f
cc_151 N_C_c_132_n N_A_c_381_n 9.00742e-19
cc_152 N_C_c_133_n N_A_c_381_n 3.9734e-19
cc_153 N_C_c_156_p N_A_c_381_n 0.00207353f
cc_154 N_C_c_161_p N_A_c_381_n 6.32429e-19
cc_155 N_C_c_156_p N_A_c_386_n 5.4333e-19
cc_156 N_C_c_133_n N_BI_c_443_n 2.41407e-19
cc_157 N_C_c_133_n N_BI_c_447_n 4.13621e-19
cc_158 N_C_c_156_p N_BI_c_450_n 6.74177e-19
cc_159 N_C_c_156_p N_BI_c_451_n 0.00240592f
cc_160 N_C_c_158_p N_B_c_563_n 0.00168372f
cc_161 N_C_c_133_n N_B_c_563_n 0.0027048f
cc_162 N_C_c_156_p N_B_c_563_n 0.00182275f
cc_163 N_C_c_161_p N_B_c_563_n 2.1095e-19
cc_164 N_C_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_165 N_C_c_158_p N_Z_XI2.X0_D 3.48267e-19
cc_166 N_C_c_178_p N_Z_XI2.X0_D 3.48267e-19
cc_167 N_C_c_132_n N_Z_XI2.X0_D 3.43419e-19
cc_168 N_C_XI3.X0_S N_Z_c_624_n 3.48267e-19
cc_169 N_C_c_158_p N_Z_c_624_n 3.41702e-19
cc_170 N_C_c_178_p N_Z_c_624_n 5.7093e-19
cc_171 N_VSS_XI9.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_172 N_VSS_c_201_n N_CI_XI10.X0_D 3.48267e-19
cc_173 N_VSS_XI7.X0_S N_CI_XI4.X0_S 3.43419e-19
cc_174 N_VSS_c_213_n N_CI_XI4.X0_S 3.48267e-19
cc_175 N_VSS_XI9.X0_S N_CI_c_316_n 3.48267e-19
cc_176 N_VSS_c_195_n N_CI_c_316_n 5.78167e-19
cc_177 N_VSS_c_201_n N_CI_c_316_n 0.00107566f
cc_178 N_VSS_c_231_n N_CI_c_316_n 0.0020072f
cc_179 N_VSS_c_233_n N_CI_c_316_n 3.32126e-19
cc_180 N_VSS_XI7.X0_S N_CI_c_334_n 3.48267e-19
cc_181 N_VSS_c_213_n N_CI_c_334_n 9.13167e-19
cc_182 N_VSS_c_205_n N_CI_c_320_n 0.00134034f
cc_183 N_VSS_c_216_n N_CI_c_320_n 0.00393483f
cc_184 N_VSS_c_235_n N_CI_c_338_n 0.00292666f
cc_185 N_VSS_c_220_n N_A_c_387_n 0.00236445f
cc_186 N_VSS_XI8.X0_PGD N_A_c_362_n 3.86211e-19
cc_187 N_VSS_XI7.X0_S N_A_c_363_n 9.18655e-19
cc_188 N_VSS_c_213_n N_A_c_363_n 0.00149545f
cc_189 N_VSS_c_216_n N_A_c_363_n 2.12774e-19
cc_190 N_VSS_c_240_n N_A_c_363_n 2.27118e-19
cc_191 N_VSS_c_205_n N_A_c_372_n 4.58305e-19
cc_192 N_VSS_c_220_n N_A_c_372_n 4.30193e-19
cc_193 N_VSS_c_287_p N_A_c_374_n 8.53264e-19
cc_194 N_VSS_c_205_n N_A_c_374_n 4.26083e-19
cc_195 N_VSS_c_220_n N_A_c_374_n 7.20776e-19
cc_196 N_VSS_XI9.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_197 N_VSS_c_201_n N_BI_XI5.X0_D 3.48267e-19
cc_198 N_VSS_XI9.X0_S N_BI_c_443_n 3.48267e-19
cc_199 N_VSS_c_201_n N_BI_c_443_n 0.00102079f
cc_200 N_VSS_c_240_n N_BI_c_443_n 3.31365e-19
cc_201 N_VSS_c_216_n N_BI_c_457_n 2.90278e-19
cc_202 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_203 N_VSS_c_213_n N_AI_XI8.X0_D 3.48267e-19
cc_204 N_VSS_XI6.X0_PGD N_AI_XI2.X0_PGD 2.84687e-19
cc_205 N_VSS_c_213_n N_AI_XI2.X0_PGD 2.04949e-19
cc_206 N_VSS_c_192_n N_AI_c_523_n 2.84687e-19
cc_207 N_VSS_XI7.X0_S N_AI_c_514_n 3.48267e-19
cc_208 N_VSS_c_205_n N_AI_c_514_n 0.00163244f
cc_209 N_VSS_c_213_n N_AI_c_514_n 0.00129029f
cc_210 N_VSS_c_213_n N_AI_c_517_n 0.00168777f
cc_211 N_VSS_c_213_n N_AI_c_528_n 2.82216e-19
cc_212 N_VSS_c_216_n N_AI_c_518_n 0.00857137f
cc_213 N_VSS_c_224_n N_B_XI6.X0_CG 0.00272012f
cc_214 N_VSS_XI8.X0_PGD N_B_c_559_n 2.07132e-19
cc_215 N_VSS_XI6.X0_PGD N_B_c_559_n 3.923e-19
cc_216 N_VSS_c_224_n N_B_c_571_n 0.00138168f
cc_217 N_VSS_c_209_n B 5.92764e-19
cc_218 N_VSS_c_224_n N_B_c_562_n 6.1245e-19
cc_219 N_VSS_c_209_n N_B_c_563_n 6.44904e-19
cc_220 N_CI_c_316_n N_BI_c_443_n 0.00104494f
cc_221 N_CI_c_324_n N_BI_c_459_n 6.86101e-19
cc_222 N_CI_c_334_n N_BI_c_447_n 8.7e-19
cc_223 N_CI_c_320_n N_BI_c_447_n 9.27611e-19
cc_224 N_CI_c_324_n N_BI_c_450_n 0.00228179f
cc_225 N_CI_c_316_n N_AI_c_514_n 5.24832e-19
cc_226 N_CI_c_334_n N_AI_c_514_n 5.10362e-19
cc_227 N_CI_c_334_n N_AI_c_517_n 0.00202744f
cc_228 N_CI_c_320_n N_AI_c_517_n 0.00654866f
cc_229 N_CI_c_324_n N_AI_c_517_n 0.00288502f
cc_230 N_CI_c_349_p N_AI_c_517_n 8.49574e-19
cc_231 N_CI_c_320_n N_AI_c_518_n 9.37419e-19
cc_232 N_CI_c_324_n N_B_c_575_n 0.00103435f
cc_233 N_CI_c_324_n N_B_c_576_n 2.42418e-19
cc_234 N_CI_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_235 N_CI_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_236 N_CI_c_334_n N_Z_XI4.X0_D 3.48267e-19
cc_237 N_CI_c_356_p N_Z_XI4.X0_D 3.48267e-19
cc_238 N_CI_XI4.X0_S N_Z_c_624_n 3.48267e-19
cc_239 N_CI_XI1.X0_S N_Z_c_624_n 3.48267e-19
cc_240 N_CI_c_334_n N_Z_c_624_n 5.68744e-19
cc_241 N_CI_c_356_p N_Z_c_624_n 5.68744e-19
cc_242 N_A_XI3.X0_PGD N_BI_XI3.X0_CG 8.79767e-19
cc_243 N_A_c_399_p N_BI_XI3.X0_CG 0.00237738f
cc_244 N_A_c_399_p N_BI_c_465_n 0.00117691f
cc_245 N_A_c_363_n N_BI_c_443_n 4.0484e-19
cc_246 N_A_c_370_n N_BI_c_443_n 6.63236e-19
cc_247 N_A_c_363_n N_BI_c_468_n 2.37396e-19
cc_248 N_A_c_386_n N_BI_c_459_n 7.92141e-19
cc_249 N_A_c_399_p N_BI_c_459_n 4.87897e-19
cc_250 N_A_c_363_n N_BI_c_471_n 3.8563e-19
cc_251 N_A_XI3.X0_PGD N_BI_c_472_n 0.00133285f
cc_252 N_A_c_386_n N_BI_c_472_n 4.79282e-19
cc_253 N_A_c_399_p N_BI_c_472_n 0.00152548f
cc_254 N_A_c_370_n N_BI_c_447_n 0.00181644f
cc_255 N_A_c_363_n N_BI_c_457_n 0.00247154f
cc_256 N_A_c_370_n N_BI_c_477_n 2.27623e-19
cc_257 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174824f
cc_258 N_A_c_370_n N_AI_XI2.X0_PGD 8.597e-19
cc_259 N_A_c_415_p N_AI_c_523_n 0.00199346f
cc_260 N_A_c_381_n N_AI_c_523_n 0.00123218f
cc_261 N_A_c_417_p N_AI_c_513_n 0.00202303f
cc_262 N_A_c_363_n N_AI_c_514_n 0.00165136f
cc_263 N_A_c_363_n N_AI_c_517_n 0.00184834f
cc_264 N_A_c_362_n N_B_c_559_n 0.00360254f
cc_265 N_A_c_363_n N_B_c_559_n 5.41329e-19
cc_266 N_A_c_374_n N_B_c_561_n 4.14098e-19
cc_267 N_A_c_381_n N_B_c_580_n 2.74862e-19
cc_268 N_A_XI3.X0_PGD N_B_c_581_n 8.79767e-19
cc_269 N_A_c_363_n B 6.972e-19
cc_270 N_A_c_370_n B 3.89684e-19
cc_271 N_A_c_370_n N_B_c_584_n 3.55503e-19
cc_272 N_A_c_381_n N_B_c_584_n 4.94081e-19
cc_273 N_A_c_381_n N_B_c_575_n 3.26384e-19
cc_274 N_A_c_362_n N_B_c_562_n 2.86506e-19
cc_275 N_A_c_370_n N_B_c_562_n 6.34732e-19
cc_276 N_A_c_370_n N_B_c_589_n 3.37713e-19
cc_277 N_A_XI3.X0_PGD N_B_c_590_n 0.00133285f
cc_278 N_A_c_370_n N_B_c_563_n 0.00206097f
cc_279 N_A_c_381_n N_B_c_563_n 0.00238641f
cc_280 N_A_c_381_n N_Z_XI2.X0_D 6.94686e-19
cc_281 N_A_XI3.X0_PGD N_Z_c_624_n 6.45939e-19
cc_282 N_A_c_370_n N_Z_c_624_n 0.00131646f
cc_283 N_A_c_381_n N_Z_c_624_n 0.00121415f
cc_284 N_BI_c_478_p N_AI_XI2.X0_PGD 8.79767e-19
cc_285 N_BI_c_471_n N_AI_XI2.X0_PGD 0.00133285f
cc_286 N_BI_c_471_n N_AI_c_546_n 6.37981e-19
cc_287 N_BI_c_457_n N_AI_c_514_n 8.05284e-19
cc_288 N_BI_c_468_n N_AI_c_517_n 4.93364e-19
cc_289 N_BI_c_447_n N_AI_c_517_n 0.00402897f
cc_290 N_BI_c_477_n N_AI_c_517_n 4.42808e-19
cc_291 N_BI_c_478_p N_AI_c_528_n 0.00234569f
cc_292 N_BI_c_468_n N_AI_c_528_n 4.6759e-19
cc_293 N_BI_c_471_n N_AI_c_528_n 0.00166302f
cc_294 N_BI_c_443_n B 4.30856e-19
cc_295 N_BI_c_447_n B 3.14738e-19
cc_296 N_BI_c_468_n N_B_c_584_n 5.92939e-19
cc_297 N_BI_c_477_n N_B_c_584_n 3.24098e-19
cc_298 N_BI_c_459_n N_B_c_575_n 0.0018551f
cc_299 N_BI_c_471_n N_B_c_589_n 0.00266367f
cc_300 N_BI_c_472_n N_B_c_589_n 6.17967e-19
cc_301 N_BI_c_471_n N_B_c_590_n 7.16621e-19
cc_302 N_BI_c_472_n N_B_c_590_n 0.00243799f
cc_303 N_BI_c_443_n N_B_c_563_n 0.00165434f
cc_304 N_BI_c_459_n N_B_c_563_n 0.00159414f
cc_305 N_BI_c_447_n N_B_c_563_n 0.0157983f
cc_306 N_BI_c_450_n N_B_c_563_n 6.88876e-19
cc_307 N_BI_c_451_n N_B_c_563_n 8.27361e-19
cc_308 N_BI_c_477_n N_B_c_607_n 0.00346365f
cc_309 N_BI_c_503_p N_B_c_607_n 0.00194674f
cc_310 N_BI_c_468_n N_B_c_576_n 3.02576e-19
cc_311 N_BI_c_450_n N_B_c_576_n 8.19447e-19
cc_312 N_BI_c_468_n N_Z_c_624_n 0.00155391f
cc_313 N_BI_c_459_n N_Z_c_624_n 0.00136914f
cc_314 N_BI_c_472_n N_Z_c_624_n 8.66889e-19
cc_315 N_BI_c_477_n N_Z_c_624_n 4.81308e-19
cc_316 N_AI_XI2.X0_PGD N_B_XI2.X0_CG 8.63152e-19
cc_317 N_AI_XI2.X0_PGD N_B_c_589_n 0.00133285f
cc_318 N_AI_XI2.X0_PGD N_Z_c_624_n 3.30612e-19
cc_319 N_B_c_584_n N_Z_c_624_n 0.00130267f
cc_320 N_B_c_575_n N_Z_c_624_n 0.00130267f
cc_321 N_B_c_589_n N_Z_c_624_n 8.66889e-19
cc_322 N_B_c_590_n N_Z_c_624_n 8.66889e-19
cc_323 N_B_c_563_n N_Z_c_624_n 0.00103251f
cc_324 N_B_c_607_n N_Z_c_624_n 0.00216955f
cc_325 N_B_c_576_n N_Z_c_624_n 9.92382e-19
*
.ends
*
*
.subckt XNOR3_HPNW1 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XNOR3_N1
.ends
*
* File: G4_XOR2_N1.pex.netlist
* Created: Fri Mar 18 15:34:38 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XOR2_N1_VSS 2 5 9 12 16 32 33 35 42 43 66 71 76 81 86 95 100 113
+ 115 116 117 122 123 128 138 140 145 146 147 150 Vss
c105 148 Vss 6.13404e-19
c106 147 Vss 3.75522e-19
c107 146 Vss 4.28045e-19
c108 145 Vss 0.0035844f
c109 140 Vss 0.00192576f
c110 138 Vss 0.00847727f
c111 128 Vss 0.00326939f
c112 123 Vss 8.39752e-19
c113 122 Vss 0.00163882f
c114 117 Vss 8.17785e-19
c115 116 Vss 0.00399757f
c116 115 Vss 0.00448448f
c117 113 Vss 0.00145652f
c118 100 Vss 0.00421853f
c119 95 Vss 0.00425358f
c120 86 Vss 1.76201e-20
c121 81 Vss 0.00164759f
c122 76 Vss 7.42069e-19
c123 71 Vss 9.70701e-19
c124 66 Vss 0.0014444f
c125 43 Vss 0.033325f
c126 42 Vss 0.0990681f
c127 35 Vss 7.82991e-20
c128 33 Vss 0.0341879f
c129 32 Vss 0.0981149f
c130 16 Vss 0.00276316f
c131 12 Vss 0.00263275f
c132 9 Vss 0.165244f
c133 5 Vss 0.166856f
c134 2 Vss 0.00267051f
r135 145 150 0.326018
r136 144 145 4.16786
r137 140 144 0.655813
r138 139 148 0.494161
r139 138 150 0.326018
r140 138 139 13.0037
r141 134 148 0.128424
r142 129 147 0.494161
r143 128 148 0.494161
r144 128 129 7.46046
r145 124 147 0.128424
r146 122 147 0.494161
r147 122 123 4.37625
r148 118 146 0.0828784
r149 116 130 0.652036
r150 116 117 10.1279
r151 115 123 0.652036
r152 114 146 0.551426
r153 114 115 12.4619
r154 113 146 0.551426
r155 112 117 0.652036
r156 112 113 4.16786
r157 86 140 1.82344
r158 81 134 4.83471
r159 76 100 1.16709
r160 76 130 2.16729
r161 71 95 1.16709
r162 71 124 2.16729
r163 66 118 1.82344
r164 45 100 0.238214
r165 43 45 1.45875
r166 42 46 0.652036
r167 42 45 1.45875
r168 39 43 0.652036
r169 35 95 0.238214
r170 33 35 1.45875
r171 32 36 0.652036
r172 32 35 1.45875
r173 29 33 0.652036
r174 16 86 1.16709
r175 12 81 1.16709
r176 9 46 2.5674
r177 9 39 2.5674
r178 5 36 2.5674
r179 5 29 2.5674
r180 2 66 1.16709
.ends

.subckt PM_G4_XOR2_N1_VDD 3 6 8 11 16 32 42 43 66 68 69 70 73 75 76 79 81 85 89
+ 91 93 98 99 100 103 109 114 Vss
c106 114 Vss 0.00542312f
c107 109 Vss 0.00583104f
c108 101 Vss 8.76285e-19
c109 100 Vss 2.39889e-19
c110 99 Vss 3.56526e-19
c111 98 Vss 0.00433275f
c112 93 Vss 0.00130328f
c113 91 Vss 0.0132502f
c114 89 Vss 0.0018632f
c115 85 Vss 7.3942e-19
c116 81 Vss 0.00447795f
c117 79 Vss 0.00129126f
c118 76 Vss 8.63329e-19
c119 75 Vss 0.00575889f
c120 73 Vss 0.00159649f
c121 70 Vss 8.67402e-19
c122 69 Vss 0.00219856f
c123 68 Vss 0.00201914f
c124 66 Vss 0.0065263f
c125 43 Vss 0.0341287f
c126 42 Vss 0.099962f
c127 33 Vss 0.0348624f
c128 32 Vss 0.0999592f
c129 16 Vss 0.00189547f
c130 11 Vss 0.165401f
c131 8 Vss 0.00162509f
c132 6 Vss 0.00218552f
c133 3 Vss 0.165774f
r134 98 103 0.349767
r135 97 98 4.16786
r136 93 103 0.306046
r137 93 95 1.82344
r138 92 101 0.494161
r139 91 97 0.652036
r140 91 92 13.0037
r141 87 101 0.128424
r142 87 89 4.83471
r143 85 114 1.16709
r144 83 85 2.16729
r145 82 100 0.494161
r146 81 101 0.494161
r147 81 82 7.46046
r148 79 109 1.16709
r149 77 100 0.128424
r150 77 79 2.16729
r151 75 83 0.652036
r152 75 76 10.1279
r153 71 99 0.0828784
r154 71 73 1.82344
r155 69 100 0.494161
r156 69 70 4.37625
r157 68 76 0.652036
r158 67 99 0.551426
r159 67 68 4.16786
r160 66 99 0.551426
r161 65 70 0.652036
r162 65 66 12.4619
r163 45 114 0.238214
r164 43 45 1.45875
r165 42 46 0.652036
r166 42 45 1.45875
r167 39 43 0.652036
r168 35 109 0.238214
r169 33 35 1.45875
r170 32 36 0.652036
r171 32 35 1.45875
r172 29 33 0.652036
r173 16 95 1.16709
r174 11 46 2.5674
r175 11 39 2.5674
r176 8 89 1.16709
r177 6 73 1.02121
r178 3 36 2.5674
r179 3 29 2.5674
.ends

.subckt PM_G4_XOR2_N1_A 2 4 7 10 18 21 24 28 39 48 54 57 62 67 72 77 85 Vss
c59 85 Vss 4.11933e-19
c60 77 Vss 9.32916e-19
c61 72 Vss 0.00720976f
c62 67 Vss 0.00368523f
c63 62 Vss 0.0024107f
c64 57 Vss 0.00389164f
c65 54 Vss 7.92361e-19
c66 48 Vss 0.126059f
c67 43 Vss 0.0296049f
c68 39 Vss 2.69463e-19
c69 28 Vss 0.152395f
c70 24 Vss 2.35358e-19
c71 21 Vss 0.169387f
c72 18 Vss 0.0715834f
c73 16 Vss 0.0247918f
c74 10 Vss 0.0674191f
c75 7 Vss 0.219218f
c76 4 Vss 0.08397f
r77 81 85 0.653045
r78 62 77 1.16709
r79 62 85 4.9014
r80 57 72 1.16709
r81 57 81 8.169
r82 51 67 1.16709
r83 51 54 0.0364688
r84 47 72 0.262036
r85 47 48 2.334
r86 44 47 2.20433
r87 39 77 0.404964
r88 33 48 0.00605528
r89 31 44 0.00605528
r90 29 43 0.494161
r91 28 30 0.652036
r92 28 29 4.84305
r93 25 43 0.128424
r94 24 67 0.0476429
r95 22 24 0.326018
r96 22 24 0.1167
r97 21 43 0.494161
r98 21 24 6.7686
r99 18 67 0.357321
r100 16 24 0.326018
r101 16 18 0.40845
r102 10 39 2.04225
r103 7 33 2.5674
r104 7 31 2.5674
r105 7 30 2.5674
r106 4 25 2.5674
r107 2 18 2.15895
.ends

.subckt PM_G4_XOR2_N1_NET1 2 7 10 31 35 44 49 58 76 Vss
c41 76 Vss 3.74063e-19
c42 58 Vss 0.00478125f
c43 49 Vss 0.00566108f
c44 44 Vss 0.0016591f
c45 35 Vss 0.102425f
c46 31 Vss 0.123619f
c47 10 Vss 0.181762f
c48 7 Vss 0.270505f
c49 2 Vss 0.00157712f
r50 72 76 0.653045
r51 49 58 1.16709
r52 49 76 12.9148
r53 44 72 2.08393
r54 33 35 1.70187
r55 30 58 0.262036
r56 30 31 2.20433
r57 27 30 2.334
r58 25 35 0.17282
r59 24 31 0.00605528
r60 21 33 0.17282
r61 18 27 0.00605528
r62 10 21 5.77665
r63 7 25 4.4346
r64 7 24 2.5674
r65 7 18 2.5674
r66 2 44 1.16709
.ends

.subckt PM_G4_XOR2_N1_NET2 2 6 9 21 22 32 33 42 47 56 74 Vss
c46 74 Vss 3.38305e-19
c47 56 Vss 0.00607606f
c48 47 Vss 0.00639628f
c49 42 Vss 0.00204719f
c50 33 Vss 0.126868f
c51 22 Vss 0.0327936f
c52 21 Vss 0.172441f
c53 9 Vss 0.361367f
c54 6 Vss 0.09048f
c55 2 Vss 0.00157712f
r56 70 74 0.660011
r57 47 56 1.16709
r58 47 74 11.3611
r59 42 70 1.95889
r60 32 56 0.262036
r61 32 33 2.26917
r62 29 32 2.26917
r63 26 33 0.00605528
r64 24 29 0.00605528
r65 21 23 0.652036
r66 21 22 4.84305
r67 18 22 0.652036
r68 9 26 2.5674
r69 9 24 2.5674
r70 9 23 7.4688
r71 6 18 2.97585
r72 2 42 1.16709
.ends

.subckt PM_G4_XOR2_N1_B 2 4 7 10 19 20 28 31 36 47 49 52 55 58 61 Vss
c39 61 Vss 0.0281877f
c40 58 Vss 0.00108886f
c41 52 Vss 0.0966253f
c42 49 Vss 0.0299431f
c43 47 Vss 0.131329f
c44 36 Vss 0.043285f
c45 31 Vss 2.35358e-19
c46 28 Vss 0.117434f
c47 20 Vss 0.03478f
c48 19 Vss 0.169387f
c49 10 Vss 0.155214f
c50 7 Vss 0.215531f
c51 4 Vss 0.0714224f
c52 2 Vss 0.083716f
r53 58 61 1.16709
r54 55 58 0.0729375
r55 50 52 2.04225
r56 45 47 4.53833
r57 40 47 0.00605528
r58 37 52 0.0685365
r59 36 50 0.0685365
r60 35 49 0.494161
r61 35 36 1.69215
r62 33 49 0.494161
r63 32 45 0.00605528
r64 31 61 0.181909
r65 29 61 0.494161
r66 29 31 0.1167
r67 28 49 0.128424
r68 28 31 4.72635
r69 23 61 0.128424
r70 23 61 0.40845
r71 22 61 0.181909
r72 20 22 6.7686
r73 19 61 0.494161
r74 19 22 0.1167
r75 16 20 0.652036
r76 10 37 5.0181
r77 7 40 2.5674
r78 7 33 2.5674
r79 7 32 2.5674
r80 4 61 2.15895
r81 2 16 2.5674
.ends

.subckt PM_G4_XOR2_N1_Z 2 4 30 33 Vss
c26 30 Vss 0.00301247f
c27 4 Vss 0.00253802f
c28 2 Vss 0.00148239f
r29 33 35 3.12589
r30 30 33 5.16814
r31 4 35 1.16709
r32 2 30 1.16709
.ends

.subckt G4_XOR2_N1  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI1.X0 N_NET1_XI1.X0_D N_VDD_XI1.X0_PGD N_B_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW1
XI9.X0 N_NET2_XI9.X0_D N_VSS_XI9.X0_PGD N_A_XI9.X0_CG N_VSS_XI9.X0_PGD
+ N_VDD_XI9.X0_S TIGFET_HPNW1
XI10.X0 N_NET1_XI1.X0_D N_VSS_XI10.X0_PGD N_B_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW1
XI3.X0 N_NET2_XI9.X0_D N_VDD_XI3.X0_PGD N_A_XI3.X0_CG N_VDD_XI3.X0_PGD
+ N_VSS_XI3.X0_S TIGFET_HPNW1
XI5.X0 N_Z_XI5.X0_D N_B_XI5.X0_PGD N_NET2_XI5.X0_CG N_B_XI5.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW1
XI8.X0 N_Z_XI8.X0_D N_A_XI8.X0_PGD N_B_XI8.X0_CG N_A_XI8.X0_PGD N_VSS_XI3.X0_S
+ TIGFET_HPNW1
XI11.X0 N_Z_XI5.X0_D N_NET1_XI11.X0_PGD N_A_XI11.X0_CG N_NET1_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW1
XI7.X0 N_Z_XI8.X0_D N_NET2_XI7.X0_PGD N_NET1_XI7.X0_CG N_NET2_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW1
*
x_PM_G4_XOR2_N1_VSS N_VSS_XI1.X0_S N_VSS_XI9.X0_PGD N_VSS_XI10.X0_PGD
+ N_VSS_XI3.X0_S N_VSS_XI7.X0_S N_VSS_c_8_p N_VSS_c_23_p N_VSS_c_56_p
+ N_VSS_c_40_p N_VSS_c_7_p N_VSS_c_3_p N_VSS_c_13_p N_VSS_c_30_p N_VSS_c_4_p
+ N_VSS_c_6_p N_VSS_c_14_p N_VSS_c_31_p N_VSS_c_10_p N_VSS_c_11_p N_VSS_c_18_p
+ N_VSS_c_19_p N_VSS_c_26_p N_VSS_c_29_p N_VSS_c_27_p N_VSS_c_62_p N_VSS_c_46_p
+ N_VSS_c_83_p N_VSS_c_12_p N_VSS_c_28_p VSS Vss PM_G4_XOR2_N1_VSS
x_PM_G4_XOR2_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI9.X0_S N_VDD_XI10.X0_S
+ N_VDD_XI3.X0_PGD N_VDD_XI11.X0_S N_VDD_c_112_n N_VDD_c_163_p N_VDD_c_113_n
+ N_VDD_c_114_n N_VDD_c_118_n N_VDD_c_121_n N_VDD_c_124_n N_VDD_c_125_n
+ N_VDD_c_127_n N_VDD_c_134_n N_VDD_c_135_n N_VDD_c_137_n N_VDD_c_141_n
+ N_VDD_c_144_n N_VDD_c_168_p N_VDD_c_149_n N_VDD_c_182_p N_VDD_c_152_n
+ N_VDD_c_153_n VDD N_VDD_c_154_n N_VDD_c_156_n Vss PM_G4_XOR2_N1_VDD
x_PM_G4_XOR2_N1_A N_A_XI9.X0_CG N_A_XI3.X0_CG N_A_XI8.X0_PGD N_A_XI11.X0_CG
+ N_A_c_212_n N_A_c_213_n N_A_c_215_n N_A_c_216_n N_A_c_246_p N_A_c_231_n A
+ N_A_c_219_n N_A_c_223_n N_A_c_224_n N_A_c_239_n N_A_c_242_p N_A_c_240_n Vss
+ PM_G4_XOR2_N1_A
x_PM_G4_XOR2_N1_NET1 N_NET1_XI1.X0_D N_NET1_XI11.X0_PGD N_NET1_XI7.X0_CG
+ N_NET1_c_282_n N_NET1_c_302_p N_NET1_c_273_n N_NET1_c_276_n N_NET1_c_289_n
+ N_NET1_c_277_n Vss PM_G4_XOR2_N1_NET1
x_PM_G4_XOR2_N1_NET2 N_NET2_XI9.X0_D N_NET2_XI5.X0_CG N_NET2_XI7.X0_PGD
+ N_NET2_c_333_n N_NET2_c_352_p N_NET2_c_334_n N_NET2_c_335_n N_NET2_c_314_n
+ N_NET2_c_318_n N_NET2_c_338_n N_NET2_c_321_n Vss PM_G4_XOR2_N1_NET2
x_PM_G4_XOR2_N1_B N_B_XI1.X0_CG N_B_XI10.X0_CG N_B_XI5.X0_PGD N_B_XI8.X0_CG
+ N_B_c_360_n N_B_c_381_n N_B_c_362_n N_B_c_363_n N_B_c_392_n N_B_c_364_n
+ N_B_c_393_n N_B_c_383_n B N_B_c_365_n N_B_c_367_n Vss PM_G4_XOR2_N1_B
x_PM_G4_XOR2_N1_Z N_Z_XI5.X0_D N_Z_XI8.X0_D N_Z_c_401_n Z Vss PM_G4_XOR2_N1_Z
cc_1 N_VSS_XI9.X0_PGD N_VDD_XI1.X0_PGD 2.77144e-19
cc_2 N_VSS_XI10.X0_PGD N_VDD_XI1.X0_PGD 0.00167677f
cc_3 N_VSS_c_3_p N_VDD_XI9.X0_S 2.05974e-19
cc_4 N_VSS_c_4_p N_VDD_XI10.X0_S 2.02468e-19
cc_5 N_VSS_XI9.X0_PGD N_VDD_XI3.X0_PGD 0.00169392f
cc_6 N_VSS_c_6_p N_VDD_XI11.X0_S 2.02468e-19
cc_7 N_VSS_c_7_p N_VDD_c_112_n 0.00167677f
cc_8 N_VSS_c_8_p N_VDD_c_113_n 0.00169392f
cc_9 N_VSS_c_3_p N_VDD_c_114_n 0.00187494f
cc_10 N_VSS_c_10_p N_VDD_c_114_n 0.00305883f
cc_11 N_VSS_c_11_p N_VDD_c_114_n 0.00593001f
cc_12 N_VSS_c_12_p N_VDD_c_114_n 8.91588e-19
cc_13 N_VSS_c_13_p N_VDD_c_118_n 4.43871e-19
cc_14 N_VSS_c_14_p N_VDD_c_118_n 3.66936e-19
cc_15 N_VSS_c_11_p N_VDD_c_118_n 0.0030181f
cc_16 N_VSS_XI1.X0_S N_VDD_c_121_n 3.7884e-19
cc_17 N_VSS_c_3_p N_VDD_c_121_n 4.73473e-19
cc_18 N_VSS_c_18_p N_VDD_c_121_n 0.00352628f
cc_19 N_VSS_c_19_p N_VDD_c_124_n 0.0010586f
cc_20 N_VSS_XI1.X0_S N_VDD_c_125_n 2.02468e-19
cc_21 N_VSS_c_3_p N_VDD_c_125_n 8.57018e-19
cc_22 N_VSS_c_8_p N_VDD_c_127_n 3.60588e-19
cc_23 N_VSS_c_23_p N_VDD_c_127_n 3.60588e-19
cc_24 N_VSS_c_13_p N_VDD_c_127_n 0.00141228f
cc_25 N_VSS_c_14_p N_VDD_c_127_n 0.00112249f
cc_26 N_VSS_c_26_p N_VDD_c_127_n 0.00343125f
cc_27 N_VSS_c_27_p N_VDD_c_127_n 0.0059942f
cc_28 N_VSS_c_28_p N_VDD_c_127_n 7.74609e-19
cc_29 N_VSS_c_29_p N_VDD_c_134_n 0.00107456f
cc_30 N_VSS_c_30_p N_VDD_c_135_n 9.22488e-19
cc_31 N_VSS_c_31_p N_VDD_c_135_n 3.82294e-19
cc_32 N_VSS_c_7_p N_VDD_c_137_n 3.60588e-19
cc_33 N_VSS_c_30_p N_VDD_c_137_n 0.00161703f
cc_34 N_VSS_c_31_p N_VDD_c_137_n 2.03837e-19
cc_35 N_VSS_c_18_p N_VDD_c_137_n 0.00605426f
cc_36 N_VSS_c_13_p N_VDD_c_141_n 9.25616e-19
cc_37 N_VSS_c_4_p N_VDD_c_141_n 9.18823e-19
cc_38 N_VSS_c_14_p N_VDD_c_141_n 3.99794e-19
cc_39 N_VSS_XI3.X0_S N_VDD_c_144_n 2.21516e-19
cc_40 N_VSS_c_40_p N_VDD_c_144_n 2.69489e-19
cc_41 N_VSS_c_30_p N_VDD_c_144_n 0.0023129f
cc_42 N_VSS_c_4_p N_VDD_c_144_n 2.43341e-19
cc_43 N_VSS_c_31_p N_VDD_c_144_n 9.55109e-19
cc_44 N_VSS_XI7.X0_S N_VDD_c_149_n 2.02468e-19
cc_45 N_VSS_c_6_p N_VDD_c_149_n 2.98086e-19
cc_46 N_VSS_c_46_p N_VDD_c_149_n 0.00130737f
cc_47 N_VSS_c_11_p N_VDD_c_152_n 9.23211e-19
cc_48 N_VSS_c_18_p N_VDD_c_153_n 0.0010761f
cc_49 N_VSS_c_30_p N_VDD_c_154_n 3.48267e-19
cc_50 N_VSS_c_31_p N_VDD_c_154_n 8.0279e-19
cc_51 N_VSS_c_13_p N_VDD_c_156_n 3.48267e-19
cc_52 N_VSS_c_14_p N_VDD_c_156_n 8.07896e-19
cc_53 N_VSS_c_14_p N_A_c_212_n 0.00234108f
cc_54 N_VSS_XI9.X0_PGD N_A_c_213_n 3.99472e-19
cc_55 N_VSS_XI10.X0_PGD N_A_c_213_n 2.20169e-19
cc_56 N_VSS_c_56_p N_A_c_215_n 9.41527e-19
cc_57 N_VSS_XI10.X0_PGD N_A_c_216_n 2.20169e-19
cc_58 N_VSS_c_13_p A 5.59945e-19
cc_59 N_VSS_c_14_p A 4.56568e-19
cc_60 N_VSS_c_4_p N_A_c_219_n 0.00506909f
cc_61 N_VSS_c_11_p N_A_c_219_n 6.18143e-19
cc_62 N_VSS_c_62_p N_A_c_219_n 0.00198136f
cc_63 N_VSS_c_46_p N_A_c_219_n 2.97351e-19
cc_64 N_VSS_c_62_p N_A_c_223_n 0.00118029f
cc_65 N_VSS_c_13_p N_A_c_224_n 4.56568e-19
cc_66 N_VSS_c_14_p N_A_c_224_n 6.1245e-19
cc_67 N_VSS_XI1.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_68 N_VSS_c_3_p N_NET1_XI1.X0_D 3.48267e-19
cc_69 N_VSS_XI1.X0_S N_NET1_c_273_n 3.48267e-19
cc_70 N_VSS_c_3_p N_NET1_c_273_n 0.00108327f
cc_71 N_VSS_c_18_p N_NET1_c_273_n 3.32126e-19
cc_72 N_VSS_c_30_p N_NET1_c_276_n 0.00167316f
cc_73 N_VSS_c_10_p N_NET1_c_277_n 3.27829e-19
cc_74 N_VSS_c_18_p N_NET1_c_277_n 6.3226e-19
cc_75 N_VSS_XI3.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_76 N_VSS_c_4_p N_NET2_XI9.X0_D 3.48267e-19
cc_77 N_VSS_XI3.X0_S N_NET2_c_314_n 3.48267e-19
cc_78 N_VSS_c_4_p N_NET2_c_314_n 0.00151106f
cc_79 N_VSS_c_11_p N_NET2_c_314_n 5.08641e-19
cc_80 N_VSS_c_27_p N_NET2_c_314_n 3.31434e-19
cc_81 N_VSS_c_4_p N_NET2_c_318_n 0.00228146f
cc_82 N_VSS_c_62_p N_NET2_c_318_n 0.00565735f
cc_83 N_VSS_c_83_p N_NET2_c_318_n 0.00115259f
cc_84 N_VSS_c_13_p N_NET2_c_321_n 5.79036e-19
cc_85 N_VSS_c_27_p N_NET2_c_321_n 0.00176418f
cc_86 N_VSS_c_31_p N_B_XI10.X0_CG 0.00234108f
cc_87 N_VSS_XI10.X0_PGD N_B_XI5.X0_PGD 0.00176522f
cc_88 N_VSS_XI9.X0_PGD N_B_c_360_n 2.20169e-19
cc_89 N_VSS_XI10.X0_PGD N_B_c_360_n 3.99472e-19
cc_90 N_VSS_XI10.X0_PGD N_B_c_362_n 4.05198e-19
cc_91 N_VSS_c_31_p N_B_c_363_n 9.49637e-19
cc_92 N_VSS_c_40_p N_B_c_364_n 0.00154836f
cc_93 N_VSS_c_30_p N_B_c_365_n 5.01474e-19
cc_94 N_VSS_c_31_p N_B_c_365_n 4.56568e-19
cc_95 N_VSS_c_30_p N_B_c_367_n 4.56568e-19
cc_96 N_VSS_c_31_p N_B_c_367_n 6.1245e-19
cc_97 N_VSS_XI3.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_98 N_VSS_XI7.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_99 N_VSS_c_4_p N_Z_XI8.X0_D 3.48267e-19
cc_100 N_VSS_c_6_p N_Z_XI8.X0_D 3.48267e-19
cc_101 N_VSS_XI3.X0_S N_Z_c_401_n 3.48267e-19
cc_102 N_VSS_XI7.X0_S N_Z_c_401_n 3.48267e-19
cc_103 N_VSS_c_4_p N_Z_c_401_n 4.94062e-19
cc_104 N_VSS_c_6_p N_Z_c_401_n 5.68744e-19
cc_105 N_VSS_c_62_p N_Z_c_401_n 3.25705e-19
cc_106 N_VDD_c_156_n N_A_XI3.X0_CG 9.28877e-19
cc_107 N_VDD_XI3.X0_PGD N_A_XI8.X0_PGD 0.00157721f
cc_108 N_VDD_XI1.X0_PGD N_A_c_213_n 2.20169e-19
cc_109 N_VDD_XI3.X0_PGD N_A_c_213_n 4.04053e-19
cc_110 N_VDD_XI3.X0_PGD N_A_c_216_n 4.05198e-19
cc_111 N_VDD_c_163_p N_A_c_231_n 0.00157721f
cc_112 N_VDD_c_114_n A 3.46645e-19
cc_113 N_VDD_c_135_n A 2.52205e-19
cc_114 N_VDD_c_141_n N_A_c_219_n 5.08705e-19
cc_115 N_VDD_c_156_n N_A_c_219_n 3.5189e-19
cc_116 N_VDD_c_168_p N_A_c_223_n 8.44396e-19
cc_117 N_VDD_c_114_n N_A_c_224_n 4.71537e-19
cc_118 N_VDD_c_154_n N_A_c_224_n 4.4222e-19
cc_119 N_VDD_c_156_n N_A_c_239_n 9.06702e-19
cc_120 N_VDD_c_168_p N_A_c_240_n 0.00102412f
cc_121 N_VDD_XI10.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_122 N_VDD_c_137_n N_NET1_XI1.X0_D 3.7884e-19
cc_123 N_VDD_c_144_n N_NET1_XI1.X0_D 3.48267e-19
cc_124 N_VDD_c_168_p N_NET1_c_282_n 8.23105e-19
cc_125 N_VDD_XI10.X0_S N_NET1_c_273_n 3.48267e-19
cc_126 N_VDD_c_137_n N_NET1_c_273_n 4.58491e-19
cc_127 N_VDD_c_144_n N_NET1_c_273_n 0.00110118f
cc_128 N_VDD_c_144_n N_NET1_c_276_n 0.00124814f
cc_129 N_VDD_c_168_p N_NET1_c_276_n 0.00341061f
cc_130 N_VDD_c_182_p N_NET1_c_276_n 8.21148e-19
cc_131 N_VDD_c_144_n N_NET1_c_289_n 2.78343e-19
cc_132 N_VDD_c_168_p N_NET1_c_289_n 0.00115624f
cc_133 N_VDD_c_182_p N_NET1_c_289_n 3.70842e-19
cc_134 N_VDD_c_135_n N_NET1_c_277_n 2.90608e-19
cc_135 N_VDD_XI9.X0_S N_NET2_XI9.X0_D 3.67949e-19
cc_136 N_VDD_c_125_n N_NET2_XI9.X0_D 3.72199e-19
cc_137 N_VDD_XI9.X0_S N_NET2_c_314_n 3.9802e-19
cc_138 N_VDD_c_125_n N_NET2_c_314_n 5.226e-19
cc_139 N_VDD_c_127_n N_NET2_c_314_n 5.01863e-19
cc_140 N_VDD_c_141_n N_NET2_c_318_n 2.9893e-19
cc_141 N_VDD_c_114_n N_B_XI1.X0_CG 3.37985e-19
cc_142 N_VDD_c_154_n N_B_XI1.X0_CG 9.28877e-19
cc_143 N_VDD_XI1.X0_PGD N_B_c_360_n 4.04053e-19
cc_144 N_VDD_XI3.X0_PGD N_B_c_360_n 2.20169e-19
cc_145 N_VDD_XI3.X0_PGD N_B_c_362_n 2.20169e-19
cc_146 N_VDD_c_144_n N_B_c_364_n 2.75901e-19
cc_147 N_VDD_c_168_p N_B_c_364_n 9.79508e-19
cc_148 N_VDD_c_141_n N_B_c_365_n 2.10322e-19
cc_149 N_VDD_c_156_n N_B_c_367_n 4.24849e-19
cc_150 N_VDD_XI10.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_151 N_VDD_XI11.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_152 N_VDD_c_144_n N_Z_XI5.X0_D 3.48267e-19
cc_153 N_VDD_c_168_p N_Z_XI5.X0_D 3.7884e-19
cc_154 N_VDD_c_149_n N_Z_XI5.X0_D 3.72199e-19
cc_155 N_VDD_XI10.X0_S N_Z_c_401_n 3.48267e-19
cc_156 N_VDD_XI11.X0_S N_Z_c_401_n 3.48267e-19
cc_157 N_VDD_c_144_n N_Z_c_401_n 7.90262e-19
cc_158 N_VDD_c_168_p N_Z_c_401_n 6.5261e-19
cc_159 N_VDD_c_149_n N_Z_c_401_n 8.53368e-19
cc_160 N_A_XI11.X0_CG N_NET1_XI11.X0_PGD 4.5346e-19
cc_161 N_A_c_242_p N_NET1_XI11.X0_PGD 0.0013363f
cc_162 N_A_c_223_n N_NET1_c_276_n 0.00121138f
cc_163 N_A_c_240_n N_NET1_c_276_n 0.00197573f
cc_164 N_A_XI11.X0_CG N_NET1_c_289_n 0.00234108f
cc_165 N_A_c_246_p N_NET1_c_289_n 0.00110158f
cc_166 N_A_c_242_p N_NET1_c_289_n 0.0014909f
cc_167 N_A_c_242_p N_NET2_XI5.X0_CG 2.18475e-19
cc_168 N_A_XI8.X0_PGD N_NET2_XI7.X0_PGD 0.00161543f
cc_169 N_A_c_216_n N_NET2_XI7.X0_PGD 3.14428e-19
cc_170 N_A_c_242_p N_NET2_XI7.X0_PGD 4.01857e-19
cc_171 N_A_XI8.X0_PGD N_NET2_c_333_n 4.60549e-19
cc_172 N_A_c_246_p N_NET2_c_334_n 2.17364e-19
cc_173 N_A_c_231_n N_NET2_c_335_n 0.00161543f
cc_174 N_A_c_219_n N_NET2_c_318_n 0.00221613f
cc_175 N_A_c_223_n N_NET2_c_318_n 7.30894e-19
cc_176 N_A_c_219_n N_NET2_c_338_n 3.44698e-19
cc_177 N_A_c_239_n N_NET2_c_338_n 9.17176e-19
cc_178 N_A_c_242_p N_NET2_c_338_n 3.34137e-19
cc_179 N_A_c_216_n N_B_XI8.X0_CG 0.003858f
cc_180 N_A_c_239_n N_B_XI8.X0_CG 0.00111269f
cc_181 N_A_c_213_n N_B_c_360_n 0.00504555f
cc_182 N_A_c_224_n N_B_c_381_n 3.67702e-19
cc_183 N_A_c_216_n N_B_c_362_n 0.00373351f
cc_184 N_A_c_216_n N_B_c_383_n 0.00215664f
cc_185 N_A_c_240_n N_B_c_365_n 2.66007e-19
cc_186 N_A_c_213_n N_B_c_367_n 4.25664e-19
cc_187 N_A_c_219_n N_Z_c_401_n 0.00323423f
cc_188 N_A_c_223_n N_Z_c_401_n 0.00319047f
cc_189 N_A_c_242_p N_Z_c_401_n 8.50872e-19
cc_190 N_NET1_c_273_n N_NET2_XI9.X0_D 2.02468e-19
cc_191 N_NET1_XI11.X0_PGD N_NET2_XI5.X0_CG 3.25363e-19
cc_192 N_NET1_c_302_p N_NET2_XI7.X0_PGD 0.00868439f
cc_193 N_NET1_XI11.X0_PGD N_NET2_c_333_n 0.00320236f
cc_194 N_NET1_XI1.X0_D N_NET2_c_314_n 2.02468e-19
cc_195 N_NET1_c_273_n N_NET2_c_314_n 3.48409e-19
cc_196 N_NET1_c_276_n N_NET2_c_318_n 0.00270459f
cc_197 N_NET1_XI7.X0_CG N_NET2_c_338_n 0.00266268f
cc_198 N_NET1_XI11.X0_PGD N_B_XI5.X0_PGD 0.00188194f
cc_199 N_NET1_XI7.X0_CG N_B_XI8.X0_CG 2.72153e-19
cc_200 N_NET1_c_282_n N_B_c_364_n 0.00165596f
cc_201 N_NET1_c_302_p N_B_c_383_n 2.72153e-19
cc_202 N_NET2_XI5.X0_CG N_B_XI5.X0_PGD 0.00233046f
cc_203 N_NET2_c_333_n N_B_XI5.X0_PGD 0.00159876f
cc_204 N_NET2_XI7.X0_PGD N_B_c_392_n 4.0517e-19
cc_205 N_NET2_c_352_p N_B_c_393_n 0.00233046f
cc_206 N_NET2_XI7.X0_PGD N_B_c_383_n 0.00313315f
cc_207 N_NET2_c_352_p N_B_c_383_n 0.00171842f
cc_208 N_NET2_XI7.X0_PGD N_Z_c_401_n 0.0012119f
cc_209 N_NET2_c_333_n N_Z_c_401_n 4.14549e-19
cc_210 N_NET2_c_318_n N_Z_c_401_n 2.62894e-19
cc_211 N_B_c_383_n N_Z_c_401_n 8.74847e-19
*
.ends
*
*
.subckt XOR2_HPNW1 A B Y VDD VSS
xgate (VSS VDD A B Y) G4_XOR2_N1
.ends
*
* File: G5_XOR3_N1.pex.netlist
* Created: Sun Apr 10 19:25:53 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XOR3_N1_VDD 2 5 9 12 14 17 34 35 44 45 54 55 77 79 80 81 84 86 90
+ 93 96 98 102 104 108 114 116 118 120 121 122 128 137 142 Vss
c124 142 Vss 0.00486824f
c125 137 Vss 0.00581297f
c126 128 Vss 0.00564406f
c127 122 Vss 0.0021675f
c128 121 Vss 2.39889e-19
c129 120 Vss 4.91069e-19
c130 119 Vss 4.36646e-19
c131 116 Vss 3.56526e-19
c132 114 Vss 0.00137025f
c133 108 Vss 8.30092e-19
c134 104 Vss 0.00588096f
c135 102 Vss 0.0013924f
c136 98 Vss 0.00493548f
c137 96 Vss 0.00124955f
c138 93 Vss 0.00253806f
c139 90 Vss 0.00359127f
c140 86 Vss 0.0066064f
c141 84 Vss 0.0015095f
c142 81 Vss 8.67096e-19
c143 80 Vss 0.0091443f
c144 79 Vss 0.00867106f
c145 77 Vss 0.00186435f
c146 55 Vss 0.0350971f
c147 54 Vss 0.099468f
c148 45 Vss 0.0346156f
c149 44 Vss 0.1003f
c150 35 Vss 0.0346129f
c151 34 Vss 0.0990563f
c152 17 Vss 0.165917f
c153 14 Vss 0.00210084f
c154 12 Vss 0.00231756f
c155 9 Vss 0.16518f
c156 5 Vss 0.165156f
c157 2 Vss 0.00208065f
r158 112 114 4.83471
r159 108 142 1.16709
r160 106 122 0.128424
r161 106 108 2.16729
r162 105 121 0.494161
r163 104 112 0.652036
r164 104 105 7.46046
r165 102 137 1.16709
r166 100 121 0.128424
r167 100 102 2.16729
r168 99 120 0.494161
r169 98 122 0.494161
r170 98 99 10.3363
r171 94 119 0.0828784
r172 94 96 2.00578
r173 93 120 0.128424
r174 92 119 0.551426
r175 92 93 3.91779
r176 90 128 1.16709
r177 88 119 0.551426
r178 88 90 5.835
r179 87 118 0.326018
r180 86 120 0.494161
r181 86 87 10.1279
r182 82 116 0.0828784
r183 82 84 1.82344
r184 80 121 0.494161
r185 80 81 15.8795
r186 79 118 0.326018
r187 78 116 0.551426
r188 78 79 13.0871
r189 77 116 0.551426
r190 76 81 0.652036
r191 76 77 4.16786
r192 57 142 0.0952857
r193 55 57 1.45875
r194 54 58 0.652036
r195 54 57 1.45875
r196 51 55 0.652036
r197 47 137 0.238214
r198 45 47 1.45875
r199 44 48 0.652036
r200 44 47 1.45875
r201 41 45 0.652036
r202 37 128 0.238214
r203 35 37 1.45875
r204 34 38 0.652036
r205 34 37 1.45875
r206 31 35 0.652036
r207 17 58 2.5674
r208 17 51 2.5674
r209 14 114 1.16709
r210 12 96 1.16709
r211 9 48 2.5674
r212 9 41 2.5674
r213 5 38 2.5674
r214 5 31 2.5674
r215 2 84 1.16709
.ends

.subckt PM_G5_XOR3_N1_C 2 4 6 8 17 20 40 43 47 52 57 62 85 87 96 97 Vss
c59 97 Vss 6.9907e-19
c60 87 Vss 0.00433475f
c61 85 Vss 0.00742725f
c62 62 Vss 0.00258068f
c63 57 Vss 0.00592074f
c64 52 Vss 0.00198267f
c65 47 Vss 7.02443e-19
c66 43 Vss 6.02755e-19
c67 40 Vss 6.7024e-19
c68 20 Vss 0.220565f
c69 17 Vss 0.0783954f
c70 15 Vss 0.0247918f
c71 8 Vss 0.00236553f
c72 4 Vss 0.0830741f
r73 88 97 0.0685365
r74 87 89 0.652036
r75 87 88 10.3363
r76 85 97 0.0685365
r77 85 96 24.7154
r78 52 89 2.16729
r79 47 62 1.16709
r80 47 97 2.08393
r81 43 57 1.16709
r82 43 96 0.531835
r83 40 43 0.0833571
r84 23 57 0.238214
r85 21 23 0.326018
r86 21 23 0.1167
r87 20 24 0.652036
r88 20 23 6.7686
r89 17 23 0.262036
r90 15 23 0.326018
r91 15 17 0.05835
r92 8 52 1.16709
r93 6 62 0.8
r94 4 24 2.5674
r95 2 17 2.50905
.ends

.subckt PM_G5_XOR3_N1_VSS 3 6 11 15 18 34 37 44 45 47 54 55 73 78 83 88 93 98
+ 107 112 121 123 124 125 130 131 136 142 153 154 155 156 Vss
c131 156 Vss 3.75522e-19
c132 155 Vss 3.87529e-19
c133 154 Vss 4.4306e-19
c134 142 Vss 0.00208493f
c135 136 Vss 0.00324551f
c136 131 Vss 8.38057e-19
c137 130 Vss 0.00579302f
c138 125 Vss 8.35119e-19
c139 124 Vss 0.00509021f
c140 123 Vss 0.00330591f
c141 121 Vss 0.00273904f
c142 112 Vss 0.00381998f
c143 107 Vss 0.00405934f
c144 98 Vss 0.00484708f
c145 93 Vss 0.00171362f
c146 88 Vss 5.59372e-19
c147 83 Vss 9.83293e-19
c148 78 Vss 0.00292041f
c149 73 Vss 0.00232164f
c150 55 Vss 0.0338093f
c151 54 Vss 0.0988897f
c152 47 Vss 7.82991e-20
c153 45 Vss 0.0347002f
c154 44 Vss 0.0989329f
c155 37 Vss 6.43685e-20
c156 35 Vss 0.0349827f
c157 34 Vss 0.1003f
c158 18 Vss 0.00259162f
c159 15 Vss 0.163916f
c160 11 Vss 0.167978f
c161 6 Vss 0.00155055f
c162 3 Vss 0.167004f
r163 148 153 1.70882
r164 143 156 0.494161
r165 142 148 0.652036
r166 142 143 7.46046
r167 138 156 0.128424
r168 137 155 0.494161
r169 136 144 0.652036
r170 136 137 7.46046
r171 132 155 0.128424
r172 130 156 0.494161
r173 130 131 15.8795
r174 126 154 0.0828784
r175 124 155 0.494161
r176 124 125 13.0037
r177 123 131 0.652036
r178 122 154 0.551426
r179 122 123 10.4196
r180 121 154 0.551426
r181 120 125 0.652036
r182 120 121 6.83529
r183 93 153 2.87582
r184 88 112 1.16709
r185 88 144 2.16729
r186 83 107 1.16709
r187 83 138 2.16729
r188 78 132 4.83471
r189 73 98 1.16709
r190 73 126 4.33978
r191 57 112 0.238214
r192 55 57 1.45875
r193 54 58 0.652036
r194 54 57 1.45875
r195 51 55 0.652036
r196 47 107 0.0952857
r197 45 47 1.45875
r198 44 48 0.652036
r199 44 47 1.45875
r200 41 45 0.652036
r201 37 98 0.238214
r202 35 37 1.45875
r203 34 38 0.652036
r204 34 37 1.45875
r205 31 35 0.652036
r206 18 93 1.16709
r207 15 58 2.5674
r208 15 51 2.5674
r209 11 48 2.5674
r210 11 41 2.5674
r211 6 78 1.16709
r212 3 38 2.5674
r213 3 31 2.5674
.ends

.subckt PM_G5_XOR3_N1_CI 2 6 8 34 39 44 79 80 82 83 84 89 Vss
c62 95 Vss 1.58755e-19
c63 89 Vss 0.00511711f
c64 84 Vss 1.26921e-19
c65 83 Vss 3.02933e-19
c66 82 Vss 0.0013099f
c67 80 Vss 4.32078e-19
c68 79 Vss 0.00369198f
c69 44 Vss 0.00182014f
c70 39 Vss 0.00109627f
c71 34 Vss 0.00267797f
c72 8 Vss 0.00276539f
c73 6 Vss 0.00212882f
c74 2 Vss 0.00154772f
r75 90 95 0.494161
r76 89 91 0.652036
r77 89 90 10.3363
r78 85 95 0.128424
r79 83 95 0.494161
r80 83 84 1.70882
r81 82 84 0.652036
r82 81 82 5.33486
r83 79 81 0.652036
r84 79 80 18.9638
r85 75 80 0.652036
r86 44 91 1.66714
r87 39 85 1.66714
r88 34 75 4.33457
r89 8 44 1.16709
r90 6 39 1.16709
r91 2 34 1.16709
.ends

.subckt PM_G5_XOR3_N1_A 2 4 7 11 21 24 45 49 51 54 55 56 58 62 63 69 74 Vss
c81 74 Vss 0.00494965f
c82 69 Vss 0.00491712f
c83 63 Vss 7.45325e-19
c84 62 Vss 6.24332e-19
c85 56 Vss 0.00115533f
c86 55 Vss 0.00958405f
c87 54 Vss 0.00423116f
c88 51 Vss 0.00507608f
c89 49 Vss 0.135015f
c90 45 Vss 0.125273f
c91 24 Vss 0.213865f
c92 21 Vss 0.0724995f
c93 19 Vss 0.0247918f
c94 7 Vss 1.00758f
c95 4 Vss 0.0850321f
r96 66 74 1.16709
r97 63 66 0.750214
r98 61 69 1.16709
r99 61 62 0.513084
r100 58 61 0.0614211
r101 55 63 0.0685365
r102 55 56 10.4613
r103 53 56 0.652036
r104 53 54 8.66914
r105 51 54 0.652036
r106 51 62 10.2113
r107 47 49 4.53833
r108 44 74 0.262036
r109 44 45 2.26917
r110 41 44 2.26917
r111 36 49 0.00605528
r112 35 45 0.00605528
r113 32 47 0.00605528
r114 31 41 0.00605528
r115 27 69 0.0952857
r116 25 27 0.326018
r117 25 27 0.1167
r118 24 28 0.652036
r119 24 27 6.7686
r120 21 27 0.3335
r121 19 27 0.326018
r122 19 21 0.2334
r123 11 36 2.5674
r124 11 32 2.5674
r125 7 11 12.837
r126 7 35 2.5674
r127 7 11 12.837
r128 7 31 2.5674
r129 4 28 2.5674
r130 2 21 2.334
.ends

.subckt PM_G5_XOR3_N1_BI 2 6 8 18 21 32 37 42 52 57 66 72 73 Vss
c61 73 Vss 1.47395e-19
c62 72 Vss 8.14419e-19
c63 66 Vss 0.00107279f
c64 57 Vss 0.00255458f
c65 52 Vss 0.00234753f
c66 42 Vss 0.00105993f
c67 37 Vss 0.001668f
c68 32 Vss 0.00236426f
c69 21 Vss 0.0573997f
c70 6 Vss 0.0573997f
c71 2 Vss 0.0015046f
r72 72 73 0.655813
r73 71 72 3.501
r74 66 71 0.655813
r75 42 57 1.16709
r76 42 73 2.00578
r77 37 52 1.16709
r78 37 77 12.0712
r79 37 66 2.00578
r80 32 49 1.16709
r81 32 77 2.08393
r82 21 57 0.50025
r83 18 52 0.50025
r84 8 21 1.80885
r85 6 18 1.80885
r86 2 49 0.1
.ends

.subckt PM_G5_XOR3_N1_AI 2 7 11 31 36 37 46 51 60 70 72 82 Vss
c55 82 Vss 2.57983e-19
c56 72 Vss 0.00283715f
c57 70 Vss 0.00386641f
c58 60 Vss 0.00539669f
c59 51 Vss 0.00147157f
c60 46 Vss 0.00243924f
c61 37 Vss 0.127837f
c62 36 Vss 6.45995e-20
c63 31 Vss 0.128147f
c64 7 Vss 0.997493f
c65 2 Vss 0.0015046f
r66 78 82 0.652036
r67 72 82 8.96089
r68 70 74 0.652036
r69 70 72 4.20954
r70 60 63 0.1
r71 51 63 1.16709
r72 51 74 1.83386
r73 46 78 4.58464
r74 36 60 0.262036
r75 36 37 2.334
r76 33 36 2.20433
r77 29 31 4.53833
r78 26 37 0.00605528
r79 25 31 0.00605528
r80 22 33 0.00605528
r81 21 29 0.00605528
r82 11 26 2.5674
r83 11 22 2.5674
r84 7 11 12.837
r85 7 25 2.5674
r86 7 11 12.837
r87 7 21 2.5674
r88 2 46 1.16709
.ends

.subckt PM_G5_XOR3_N1_B 2 4 6 8 16 17 24 26 33 38 42 45 50 55 60 65 73 74 80 86
+ 91 92 Vss
c91 92 Vss 1.10364e-19
c92 91 Vss 9.61135e-19
c93 86 Vss 5.98353e-19
c94 80 Vss 8.23772e-19
c95 74 Vss 5.75465e-19
c96 73 Vss 0.00321909f
c97 65 Vss 0.00250661f
c98 60 Vss 0.00207758f
c99 55 Vss 0.00386058f
c100 50 Vss 0.00113661f
c101 45 Vss 4.31637e-19
c102 42 Vss 4.09773e-19
c103 38 Vss 5.37175e-19
c104 33 Vss 6.95992e-20
c105 26 Vss 0.0573997f
c106 24 Vss 7.82991e-20
c107 20 Vss 0.0247918f
c108 17 Vss 0.0338376f
c109 16 Vss 0.183114f
c110 8 Vss 0.0573997f
c111 4 Vss 0.0714013f
c112 2 Vss 0.0826046f
r113 90 92 0.65228
r114 90 91 3.46076
r115 86 91 0.65228
r116 73 80 0.0685365
r117 73 74 10.3363
r118 69 74 0.652036
r119 50 65 1.16709
r120 50 92 2.1395
r121 45 60 1.16709
r122 45 86 2.1006
r123 45 80 2.08393
r124 38 55 1.16709
r125 38 69 2.16729
r126 38 42 0.0729375
r127 36 55 0.0476429
r128 33 65 0.50025
r129 26 60 0.50025
r130 24 55 0.357321
r131 20 36 0.326018
r132 20 24 0.40845
r133 17 36 6.7686
r134 16 36 0.326018
r135 16 36 0.1167
r136 13 17 0.652036
r137 8 33 1.80885
r138 6 26 1.80885
r139 4 24 2.15895
r140 2 13 2.5674
.ends

.subckt PM_G5_XOR3_N1_Z 2 4 30 33 Vss
c30 30 Vss 0.00324462f
c31 4 Vss 0.00153036f
c32 2 Vss 0.00166246f
r33 33 35 4.50129
r34 30 33 4.668
r35 4 35 1.16709
r36 2 30 1.16709
.ends

.subckt G5_XOR3_N1  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI10.X0 N_CI_XI10.X0_D N_VSS_XI10.X0_PGD N_C_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW1
XI9.X0 N_CI_XI10.X0_D N_VDD_XI9.X0_PGD N_C_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW1
XI5.X0 N_BI_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW1
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW1
XI6.X0 N_BI_XI5.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW1
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW1
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_BI_XI2.X0_CG N_AI_XI2.X0_PGD N_C_XI2.X0_S
+ TIGFET_HPNW1
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_B_XI4.X0_CG N_AI_XI4.X0_PGD N_CI_XI4.X0_S
+ TIGFET_HPNW1
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_B_XI3.X0_CG N_A_XI3.X0_PGD N_C_XI3.X0_S
+ TIGFET_HPNW1
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_BI_XI1.X0_CG N_A_XI1.X0_PGD N_CI_XI1.X0_S
+ TIGFET_HPNW1
*
x_PM_G5_XOR3_N1_VDD N_VDD_XI10.X0_S N_VDD_XI9.X0_PGD N_VDD_XI5.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI6.X0_S N_VDD_XI7.X0_PGD N_VDD_c_121_p N_VDD_c_20_p
+ N_VDD_c_25_p N_VDD_c_4_p N_VDD_c_109_p N_VDD_c_21_p N_VDD_c_6_p N_VDD_c_27_p
+ N_VDD_c_5_p N_VDD_c_64_p N_VDD_c_29_p N_VDD_c_30_p N_VDD_c_31_p N_VDD_c_37_p
+ N_VDD_c_34_p N_VDD_c_22_p N_VDD_c_11_p N_VDD_c_26_p N_VDD_c_39_p N_VDD_c_12_p
+ N_VDD_c_60_p VDD N_VDD_c_68_p N_VDD_c_72_p N_VDD_c_19_p N_VDD_c_2_p
+ N_VDD_c_44_p N_VDD_c_40_p Vss PM_G5_XOR3_N1_VDD
x_PM_G5_XOR3_N1_C N_C_XI10.X0_CG N_C_XI9.X0_CG N_C_XI2.X0_S N_C_XI3.X0_S
+ N_C_c_144_p N_C_c_127_n C N_C_c_140_p N_C_c_157_p N_C_c_179_p N_C_c_132_n
+ N_C_c_134_n N_C_c_135_n N_C_c_156_p N_C_c_141_p N_C_c_160_p Vss
+ PM_G5_XOR3_N1_C
x_PM_G5_XOR3_N1_VSS N_VSS_XI10.X0_PGD N_VSS_XI9.X0_S N_VSS_XI8.X0_PGD
+ N_VSS_XI6.X0_PGD N_VSS_XI7.X0_S N_VSS_c_191_n N_VSS_c_250_n N_VSS_c_192_n
+ N_VSS_c_194_n N_VSS_c_288_p N_VSS_c_195_n N_VSS_c_196_n N_VSS_c_198_n
+ N_VSS_c_204_n N_VSS_c_208_n N_VSS_c_212_n N_VSS_c_216_n N_VSS_c_218_n
+ N_VSS_c_221_n N_VSS_c_225_n N_VSS_c_229_n N_VSS_c_232_n N_VSS_c_234_n
+ N_VSS_c_235_n N_VSS_c_236_n N_VSS_c_240_n N_VSS_c_241_n N_VSS_c_244_n VSS
+ N_VSS_c_246_n N_VSS_c_247_n N_VSS_c_248_n Vss PM_G5_XOR3_N1_VSS
x_PM_G5_XOR3_N1_CI N_CI_XI10.X0_D N_CI_XI4.X0_S N_CI_XI1.X0_S N_CI_c_317_n
+ N_CI_c_333_n N_CI_c_373_p N_CI_c_321_n N_CI_c_337_n N_CI_c_339_n N_CI_c_347_p
+ N_CI_c_356_p N_CI_c_325_n Vss PM_G5_XOR3_N1_CI
x_PM_G5_XOR3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI3.X0_PGD N_A_XI1.X0_PGD
+ N_A_c_402_n N_A_c_378_n N_A_c_428_p N_A_c_430_p N_A_c_379_n N_A_c_387_n
+ N_A_c_396_n N_A_c_388_n A N_A_c_389_n N_A_c_401_n N_A_c_390_n N_A_c_434_p Vss
+ PM_G5_XOR3_N1_A
x_PM_G5_XOR3_N1_BI N_BI_XI5.X0_D N_BI_XI2.X0_CG N_BI_XI1.X0_CG N_BI_c_480_n
+ N_BI_c_481_n N_BI_c_460_n N_BI_c_464_n N_BI_c_478_n N_BI_c_486_n N_BI_c_487_n
+ N_BI_c_467_n N_BI_c_506_p N_BI_c_479_n Vss PM_G5_XOR3_N1_BI
x_PM_G5_XOR3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_532_n
+ N_AI_c_566_p N_AI_c_522_n N_AI_c_523_n N_AI_c_537_n N_AI_c_527_n N_AI_c_528_n
+ N_AI_c_529_n N_AI_c_540_n Vss PM_G5_XOR3_N1_AI
x_PM_G5_XOR3_N1_B N_B_XI5.X0_CG N_B_XI6.X0_CG N_B_XI4.X0_CG N_B_XI3.X0_CG
+ N_B_c_576_n N_B_c_578_n N_B_c_590_n N_B_c_648_n N_B_c_611_n N_B_c_579_n B
+ N_B_c_615_n N_B_c_583_n N_B_c_580_n N_B_c_620_n N_B_c_621_n N_B_c_581_n
+ N_B_c_602_n N_B_c_603_n N_B_c_585_n N_B_c_645_n N_B_c_586_n Vss
+ PM_G5_XOR3_N1_B
x_PM_G5_XOR3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_669_n Z Vss PM_G5_XOR3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_C_XI9.X0_CG 9.6041e-19
cc_2 N_VDD_c_2_p N_C_XI9.X0_CG 8.03148e-19
cc_3 N_VDD_XI9.X0_PGD N_C_c_127_n 4.16623e-19
cc_4 N_VDD_c_4_p N_C_c_127_n 9.6041e-19
cc_5 N_VDD_c_5_p N_C_c_127_n 0.00125128f
cc_6 N_VDD_c_6_p C 4.36744e-19
cc_7 N_VDD_c_5_p C 0.00161703f
cc_8 N_VDD_c_6_p N_C_c_132_n 3.66936e-19
cc_9 N_VDD_c_5_p N_C_c_132_n 2.84956e-19
cc_10 N_VDD_XI6.X0_S N_C_c_134_n 3.43419e-19
cc_11 N_VDD_c_11_p N_C_c_135_n 4.67477e-19
cc_12 N_VDD_c_12_p N_C_c_135_n 7.7658e-19
cc_13 N_VDD_XI9.X0_PGD N_VSS_XI10.X0_PGD 0.00173038f
cc_14 N_VDD_c_5_p N_VSS_XI9.X0_S 3.7884e-19
cc_15 N_VDD_XI5.X0_PGD N_VSS_XI8.X0_PGD 2.27468e-19
cc_16 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172148f
cc_17 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017188f
cc_18 N_VDD_XI7.X0_PGD N_VSS_XI6.X0_PGD 2.1536e-19
cc_19 N_VDD_c_19_p N_VSS_XI7.X0_S 4.04413e-19
cc_20 N_VDD_c_20_p N_VSS_c_191_n 0.00173038f
cc_21 N_VDD_c_21_p N_VSS_c_192_n 0.00172148f
cc_22 N_VDD_c_22_p N_VSS_c_192_n 2.51785e-19
cc_23 N_VDD_c_22_p N_VSS_c_194_n 3.71017e-19
cc_24 N_VDD_c_12_p N_VSS_c_195_n 2.35445e-19
cc_25 N_VDD_c_25_p N_VSS_c_196_n 0.0017188f
cc_26 N_VDD_c_26_p N_VSS_c_196_n 2.74208e-19
cc_27 N_VDD_c_27_p N_VSS_c_198_n 4.32468e-19
cc_28 N_VDD_c_5_p N_VSS_c_198_n 4.60511e-19
cc_29 N_VDD_c_29_p N_VSS_c_198_n 0.00130521f
cc_30 N_VDD_c_30_p N_VSS_c_198_n 4.5978e-19
cc_31 N_VDD_c_31_p N_VSS_c_198_n 3.98949e-19
cc_32 N_VDD_c_2_p N_VSS_c_198_n 3.48267e-19
cc_33 N_VDD_c_5_p N_VSS_c_204_n 4.58491e-19
cc_34 N_VDD_c_34_p N_VSS_c_204_n 2.25587e-19
cc_35 N_VDD_c_11_p N_VSS_c_204_n 7.77634e-19
cc_36 N_VDD_c_12_p N_VSS_c_204_n 3.28649e-19
cc_37 N_VDD_c_37_p N_VSS_c_208_n 4.0876e-19
cc_38 N_VDD_c_22_p N_VSS_c_208_n 0.00141228f
cc_39 N_VDD_c_39_p N_VSS_c_208_n 8.73606e-19
cc_40 N_VDD_c_40_p N_VSS_c_208_n 3.48267e-19
cc_41 N_VDD_c_11_p N_VSS_c_212_n 6.87451e-19
cc_42 N_VDD_c_26_p N_VSS_c_212_n 0.00141228f
cc_43 N_VDD_c_12_p N_VSS_c_212_n 0.00254823f
cc_44 N_VDD_c_44_p N_VSS_c_212_n 3.48267e-19
cc_45 N_VDD_c_39_p N_VSS_c_216_n 7.30795e-19
cc_46 N_VDD_c_19_p N_VSS_c_216_n 5.00098e-19
cc_47 N_VDD_c_27_p N_VSS_c_218_n 4.41003e-19
cc_48 N_VDD_c_31_p N_VSS_c_218_n 3.89161e-19
cc_49 N_VDD_c_2_p N_VSS_c_218_n 7.99831e-19
cc_50 N_VDD_c_37_p N_VSS_c_221_n 3.48267e-19
cc_51 N_VDD_c_22_p N_VSS_c_221_n 0.00112249f
cc_52 N_VDD_c_39_p N_VSS_c_221_n 3.99794e-19
cc_53 N_VDD_c_40_p N_VSS_c_221_n 8.07559e-19
cc_54 N_VDD_c_11_p N_VSS_c_225_n 3.82294e-19
cc_55 N_VDD_c_26_p N_VSS_c_225_n 0.00112249f
cc_56 N_VDD_c_12_p N_VSS_c_225_n 9.55109e-19
cc_57 N_VDD_c_44_p N_VSS_c_225_n 8.01441e-19
cc_58 N_VDD_c_6_p N_VSS_c_229_n 0.003116f
cc_59 N_VDD_c_27_p N_VSS_c_229_n 7.60301e-19
cc_60 N_VDD_c_60_p N_VSS_c_229_n 0.0010705f
cc_61 N_VDD_c_27_p N_VSS_c_232_n 0.00754268f
cc_62 N_VDD_c_31_p N_VSS_c_232_n 9.72927e-19
cc_63 N_VDD_c_5_p N_VSS_c_234_n 0.00967241f
cc_64 N_VDD_c_64_p N_VSS_c_235_n 0.00107121f
cc_65 N_VDD_c_30_p N_VSS_c_236_n 0.0081111f
cc_66 N_VDD_c_34_p N_VSS_c_236_n 7.52646e-19
cc_67 N_VDD_c_22_p N_VSS_c_236_n 0.00375883f
cc_68 N_VDD_c_68_p N_VSS_c_236_n 0.0014027f
cc_69 N_VDD_c_27_p N_VSS_c_240_n 0.00107333f
cc_70 N_VDD_c_5_p N_VSS_c_241_n 0.00142828f
cc_71 N_VDD_c_26_p N_VSS_c_241_n 0.00543165f
cc_72 N_VDD_c_72_p N_VSS_c_241_n 0.00106247f
cc_73 N_VDD_c_22_p N_VSS_c_244_n 0.00372698f
cc_74 N_VDD_c_19_p N_VSS_c_244_n 0.00347642f
cc_75 N_VDD_c_27_p N_VSS_c_246_n 0.00112682f
cc_76 N_VDD_c_5_p N_VSS_c_247_n 0.00104966f
cc_77 N_VDD_c_22_p N_VSS_c_248_n 7.74609e-19
cc_78 N_VDD_XI10.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_79 N_VDD_c_29_p N_CI_XI10.X0_D 3.72199e-19
cc_80 N_VDD_XI10.X0_S N_CI_c_317_n 3.48267e-19
cc_81 N_VDD_c_5_p N_CI_c_317_n 5.01863e-19
cc_82 N_VDD_c_29_p N_CI_c_317_n 5.226e-19
cc_83 N_VDD_c_31_p N_CI_c_317_n 4.13481e-19
cc_84 N_VDD_c_31_p N_CI_c_321_n 7.11597e-19
cc_85 N_VDD_c_34_p N_CI_c_321_n 7.78475e-19
cc_86 N_VDD_c_40_p N_A_XI7.X0_CG 0.00119068f
cc_87 N_VDD_XI7.X0_PGD N_A_c_378_n 3.90714e-19
cc_88 N_VDD_XI6.X0_S N_A_c_379_n 2.96819e-19
cc_89 N_VDD_XI7.X0_PGD N_A_c_379_n 2.39692e-19
cc_90 N_VDD_c_22_p N_A_c_379_n 5.16693e-19
cc_91 N_VDD_c_26_p N_A_c_379_n 4.57585e-19
cc_92 N_VDD_c_39_p N_A_c_379_n 5.97577e-19
cc_93 N_VDD_c_12_p N_A_c_379_n 4.47961e-19
cc_94 N_VDD_c_19_p N_A_c_379_n 4.69788e-19
cc_95 N_VDD_c_40_p N_A_c_379_n 4.46731e-19
cc_96 N_VDD_XI6.X0_S N_A_c_387_n 9.18655e-19
cc_97 N_VDD_c_12_p N_A_c_388_n 0.00610545f
cc_98 N_VDD_c_31_p N_A_c_389_n 8.33062e-19
cc_99 N_VDD_c_31_p N_A_c_390_n 6.30148e-19
cc_100 N_VDD_c_44_p N_A_c_390_n 5.39283e-19
cc_101 N_VDD_XI6.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_102 N_VDD_c_12_p N_BI_XI5.X0_D 3.48267e-19
cc_103 N_VDD_XI6.X0_S N_BI_c_460_n 3.48267e-19
cc_104 N_VDD_c_26_p N_BI_c_460_n 4.87462e-19
cc_105 N_VDD_c_12_p N_BI_c_460_n 5.0516e-19
cc_106 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_107 N_VDD_c_22_p N_AI_XI8.X0_D 4.04413e-19
cc_108 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.98495e-19
cc_109 N_VDD_c_109_p N_AI_c_522_n 2.98495e-19
cc_110 N_VDD_XI8.X0_S N_AI_c_523_n 3.48267e-19
cc_111 N_VDD_c_34_p N_AI_c_523_n 4.96286e-19
cc_112 N_VDD_c_22_p N_AI_c_523_n 4.84258e-19
cc_113 N_VDD_c_39_p N_AI_c_523_n 5.74209e-19
cc_114 N_VDD_c_39_p N_AI_c_527_n 2.15672e-19
cc_115 N_VDD_c_19_p N_AI_c_528_n 3.25291e-19
cc_116 N_VDD_c_22_p N_AI_c_529_n 2.81017e-19
cc_117 N_VDD_XI9.X0_PGD N_B_XI5.X0_CG 9.57243e-19
cc_118 N_VDD_c_44_p N_B_XI5.X0_CG 9.74645e-19
cc_119 N_VDD_XI5.X0_PGD N_B_c_576_n 3.9688e-19
cc_120 N_VDD_XI7.X0_PGD N_B_c_576_n 2.07132e-19
cc_121 N_VDD_c_121_p N_B_c_578_n 9.57243e-19
cc_122 N_VDD_c_31_p N_B_c_579_n 6.08224e-19
cc_123 N_VDD_c_40_p N_B_c_580_n 3.47237e-19
cc_124 N_VDD_c_12_p N_B_c_581_n 2.72308e-19
cc_125 N_C_c_127_n N_VSS_XI10.X0_PGD 4.16623e-19
cc_126 N_C_c_132_n N_VSS_c_250_n 6.87259e-19
cc_127 C N_VSS_c_198_n 4.80408e-19
cc_128 N_C_c_140_p N_VSS_c_198_n 3.9981e-19
cc_129 N_C_c_141_p N_VSS_c_198_n 2.54015e-19
cc_130 N_C_c_135_n N_VSS_c_204_n 0.00185659f
cc_131 N_C_c_135_n N_VSS_c_212_n 0.00161389f
cc_132 N_C_c_144_p N_VSS_c_218_n 0.0041277f
cc_133 C N_VSS_c_218_n 4.20453e-19
cc_134 N_C_c_132_n N_VSS_c_218_n 0.00184261f
cc_135 N_C_c_140_p N_VSS_c_229_n 4.01014e-19
cc_136 N_C_c_141_p N_VSS_c_229_n 2.65147e-19
cc_137 C N_VSS_c_234_n 3.52403e-19
cc_138 N_C_c_140_p N_VSS_c_234_n 0.00136475f
cc_139 N_C_c_135_n N_VSS_c_234_n 0.00239048f
cc_140 N_C_c_141_p N_VSS_c_234_n 5.40072e-19
cc_141 N_C_c_135_n N_VSS_c_241_n 0.00182168f
cc_142 N_C_c_135_n N_CI_c_317_n 0.00135409f
cc_143 N_C_c_135_n N_CI_c_321_n 0.0042263f
cc_144 N_C_c_156_p N_CI_c_325_n 6.92841e-19
cc_145 N_C_c_157_p N_A_c_387_n 0.00149093f
cc_146 N_C_c_134_n N_A_c_387_n 8.20481e-19
cc_147 N_C_c_135_n N_A_c_387_n 2.83242e-19
cc_148 N_C_c_160_p N_A_c_387_n 2.26175e-19
cc_149 N_C_c_157_p N_A_c_396_n 0.00194268f
cc_150 N_C_c_134_n N_A_c_396_n 9.18655e-19
cc_151 N_C_c_135_n N_A_c_396_n 4.77334e-19
cc_152 N_C_c_156_p N_A_c_396_n 0.00211066f
cc_153 N_C_c_160_p N_A_c_396_n 6.30333e-19
cc_154 N_C_c_156_p N_A_c_401_n 5.46695e-19
cc_155 N_C_c_135_n N_BI_c_460_n 0.00227671f
cc_156 N_C_c_135_n N_BI_c_464_n 0.00490342f
cc_157 N_C_c_156_p N_BI_c_464_n 0.0015987f
cc_158 N_C_c_160_p N_BI_c_464_n 0.0013513f
cc_159 N_C_c_156_p N_BI_c_467_n 9.86034e-19
cc_160 N_C_c_135_n N_B_c_579_n 2.53746e-19
cc_161 N_C_c_156_p N_B_c_583_n 2.11999e-19
cc_162 N_C_c_157_p N_B_c_581_n 4.78342e-19
cc_163 N_C_c_156_p N_B_c_585_n 5.08651e-19
cc_164 N_C_c_156_p N_B_c_586_n 0.00239488f
cc_165 N_C_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_166 N_C_c_157_p N_Z_XI2.X0_D 3.48267e-19
cc_167 N_C_c_179_p N_Z_XI2.X0_D 3.48267e-19
cc_168 N_C_c_134_n N_Z_XI2.X0_D 3.43419e-19
cc_169 N_C_XI3.X0_S N_Z_c_669_n 3.48267e-19
cc_170 N_C_c_157_p N_Z_c_669_n 3.23828e-19
cc_171 N_C_c_179_p N_Z_c_669_n 5.71075e-19
cc_172 N_VSS_XI9.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_173 N_VSS_c_204_n N_CI_XI10.X0_D 3.48267e-19
cc_174 N_VSS_XI7.X0_S N_CI_XI4.X0_S 3.43419e-19
cc_175 N_VSS_c_216_n N_CI_XI4.X0_S 3.48267e-19
cc_176 N_VSS_c_198_n N_CI_c_317_n 5.88914e-19
cc_177 N_VSS_c_204_n N_CI_c_317_n 8.48865e-19
cc_178 N_VSS_c_234_n N_CI_c_317_n 3.32126e-19
cc_179 N_VSS_XI7.X0_S N_CI_c_333_n 3.48267e-19
cc_180 N_VSS_c_216_n N_CI_c_333_n 7.99744e-19
cc_181 N_VSS_c_208_n N_CI_c_321_n 3.41088e-19
cc_182 N_VSS_c_244_n N_CI_c_321_n 4.44969e-19
cc_183 N_VSS_c_232_n N_CI_c_337_n 2.78598e-19
cc_184 N_VSS_c_236_n N_CI_c_337_n 0.00159458f
cc_185 N_VSS_c_216_n N_CI_c_339_n 0.00104291f
cc_186 N_VSS_c_221_n N_A_c_402_n 0.00297797f
cc_187 N_VSS_XI8.X0_PGD N_A_c_378_n 3.85826e-19
cc_188 N_VSS_XI7.X0_S N_A_c_379_n 9.18655e-19
cc_189 N_VSS_c_216_n N_A_c_379_n 0.00131738f
cc_190 N_VSS_c_241_n N_A_c_379_n 3.01443e-19
cc_191 N_VSS_c_244_n N_A_c_379_n 5.02211e-19
cc_192 N_VSS_c_208_n N_A_c_389_n 5.62647e-19
cc_193 N_VSS_c_221_n N_A_c_389_n 4.60973e-19
cc_194 N_VSS_c_288_p N_A_c_390_n 9.36847e-19
cc_195 N_VSS_c_208_n N_A_c_390_n 4.56568e-19
cc_196 N_VSS_c_221_n N_A_c_390_n 8.15819e-19
cc_197 N_VSS_XI9.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_198 N_VSS_XI9.X0_S N_BI_c_460_n 3.48267e-19
cc_199 N_VSS_c_204_n N_BI_c_460_n 7.98486e-19
cc_200 N_VSS_c_241_n N_BI_c_460_n 3.20743e-19
cc_201 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_202 N_VSS_XI6.X0_PGD N_AI_XI2.X0_PGD 2.8463e-19
cc_203 N_VSS_c_195_n N_AI_c_532_n 2.8463e-19
cc_204 N_VSS_XI7.X0_S N_AI_c_523_n 3.48267e-19
cc_205 N_VSS_c_208_n N_AI_c_523_n 0.00108072f
cc_206 N_VSS_c_216_n N_AI_c_523_n 0.00193557f
cc_207 N_VSS_c_244_n N_AI_c_523_n 3.6914e-19
cc_208 N_VSS_c_216_n N_AI_c_537_n 8.20606e-19
cc_209 N_VSS_c_244_n N_AI_c_528_n 9.54335e-19
cc_210 N_VSS_c_244_n N_AI_c_529_n 0.00515467f
cc_211 N_VSS_c_244_n N_AI_c_540_n 0.00185629f
cc_212 N_VSS_c_225_n N_B_XI6.X0_CG 0.00272012f
cc_213 N_VSS_XI8.X0_PGD N_B_c_576_n 2.07132e-19
cc_214 N_VSS_XI6.X0_PGD N_B_c_576_n 3.923e-19
cc_215 N_VSS_c_225_n N_B_c_590_n 0.00130195f
cc_216 N_VSS_c_212_n N_B_c_579_n 7.62066e-19
cc_217 N_VSS_c_212_n B 5.66975e-19
cc_218 N_VSS_c_225_n B 4.56568e-19
cc_219 N_VSS_c_225_n N_B_c_580_n 6.1245e-19
cc_220 N_VSS_c_216_n N_B_c_581_n 6.79536e-19
cc_221 N_CI_c_339_n N_A_c_379_n 6.20926e-19
cc_222 N_CI_c_321_n N_A_c_389_n 0.00116415f
cc_223 N_CI_c_339_n N_A_c_389_n 2.08707e-19
cc_224 N_CI_c_317_n N_BI_c_460_n 5.94242e-19
cc_225 N_CI_c_321_n N_BI_c_460_n 0.00302092f
cc_226 N_CI_c_333_n N_BI_c_464_n 3.50977e-19
cc_227 N_CI_c_321_n N_BI_c_464_n 0.00752744f
cc_228 N_CI_c_347_p N_BI_c_464_n 4.80593e-19
cc_229 N_CI_c_325_n N_BI_c_464_n 5.67893e-19
cc_230 N_CI_c_325_n N_BI_c_478_n 0.00102574f
cc_231 N_CI_c_325_n N_BI_c_479_n 2.55507e-19
cc_232 N_CI_c_321_n N_AI_c_523_n 8.44506e-19
cc_233 N_CI_c_339_n N_AI_c_523_n 0.00100365f
cc_234 N_CI_c_325_n N_AI_c_537_n 0.00169084f
cc_235 N_CI_c_333_n N_AI_c_528_n 8.33462e-19
cc_236 N_CI_c_347_p N_AI_c_528_n 7.14401e-19
cc_237 N_CI_c_356_p N_AI_c_528_n 2.16882e-19
cc_238 N_CI_c_325_n N_AI_c_528_n 5.16616e-19
cc_239 N_CI_c_321_n N_AI_c_529_n 0.00115159f
cc_240 N_CI_c_356_p N_AI_c_529_n 0.00241787f
cc_241 N_CI_c_317_n N_B_c_579_n 2.7112e-19
cc_242 N_CI_c_325_n N_B_c_583_n 7.18914e-19
cc_243 N_CI_c_333_n N_B_c_581_n 8.80932e-19
cc_244 N_CI_c_321_n N_B_c_581_n 0.00348609f
cc_245 N_CI_c_347_p N_B_c_581_n 2.27019e-19
cc_246 N_CI_c_325_n N_B_c_581_n 2.27123e-19
cc_247 N_CI_c_321_n N_B_c_602_n 0.00142048f
cc_248 N_CI_c_339_n N_B_c_603_n 3.62522e-19
cc_249 N_CI_c_339_n N_B_c_585_n 4.56062e-19
cc_250 N_CI_c_325_n N_B_c_585_n 0.00270237f
cc_251 N_CI_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_252 N_CI_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_253 N_CI_c_333_n N_Z_XI4.X0_D 3.48267e-19
cc_254 N_CI_c_373_p N_Z_XI4.X0_D 3.48267e-19
cc_255 N_CI_XI4.X0_S N_Z_c_669_n 3.48267e-19
cc_256 N_CI_c_333_n N_Z_c_669_n 5.68744e-19
cc_257 N_CI_c_373_p N_Z_c_669_n 6.06579e-19
cc_258 N_A_c_396_n N_BI_c_480_n 3.17089e-19
cc_259 N_A_XI3.X0_PGD N_BI_c_481_n 8.79767e-19
cc_260 N_A_c_379_n N_BI_c_460_n 4.32688e-19
cc_261 N_A_c_387_n N_BI_c_464_n 9.32646e-19
cc_262 N_A_c_396_n N_BI_c_464_n 5.00869e-19
cc_263 N_A_c_396_n N_BI_c_478_n 3.33012e-19
cc_264 N_A_c_387_n N_BI_c_486_n 3.37713e-19
cc_265 N_A_XI3.X0_PGD N_BI_c_487_n 0.00133285f
cc_266 N_A_c_396_n N_BI_c_467_n 0.00106538f
cc_267 N_A_c_379_n N_AI_XI8.X0_D 9.18655e-19
cc_268 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174819f
cc_269 N_A_c_387_n N_AI_XI2.X0_PGD 8.52417e-19
cc_270 N_A_c_428_p N_AI_c_532_n 0.00199595f
cc_271 N_A_c_396_n N_AI_c_532_n 0.00123184f
cc_272 N_A_c_430_p N_AI_c_522_n 0.00202022f
cc_273 N_A_c_379_n N_AI_c_523_n 0.00136181f
cc_274 N_A_c_379_n N_AI_c_529_n 2.67536e-19
cc_275 N_A_XI3.X0_PGD N_B_XI3.X0_CG 8.79767e-19
cc_276 N_A_c_434_p N_B_XI3.X0_CG 0.00237738f
cc_277 N_A_c_378_n N_B_c_576_n 0.0036024f
cc_278 N_A_c_379_n N_B_c_576_n 5.40888e-19
cc_279 N_A_c_390_n N_B_c_578_n 4.08399e-19
cc_280 N_A_c_434_p N_B_c_611_n 0.00115102f
cc_281 N_A_c_387_n N_B_c_579_n 6.16253e-19
cc_282 N_A_c_379_n B 7.07944e-19
cc_283 N_A_c_387_n B 5.00495e-19
cc_284 N_A_c_379_n N_B_c_615_n 2.41829e-19
cc_285 N_A_c_401_n N_B_c_583_n 8.44727e-19
cc_286 N_A_c_434_p N_B_c_583_n 4.84491e-19
cc_287 N_A_c_378_n N_B_c_580_n 2.87365e-19
cc_288 N_A_c_387_n N_B_c_580_n 6.85754e-19
cc_289 N_A_c_379_n N_B_c_620_n 3.8563e-19
cc_290 N_A_XI3.X0_PGD N_B_c_621_n 0.00133285f
cc_291 N_A_c_401_n N_B_c_621_n 4.67029e-19
cc_292 N_A_c_434_p N_B_c_621_n 0.0014909f
cc_293 N_A_c_387_n N_B_c_581_n 0.00225059f
cc_294 N_A_c_396_n N_B_c_581_n 8.88958e-19
cc_295 N_A_c_379_n N_B_c_602_n 0.00244205f
cc_296 N_A_c_396_n N_Z_XI2.X0_D 6.94686e-19
cc_297 N_A_XI3.X0_PGD N_Z_c_669_n 6.30408e-19
cc_298 N_A_c_387_n N_Z_c_669_n 0.00124827f
cc_299 N_A_c_396_n N_Z_c_669_n 0.00121415f
cc_300 N_BI_XI2.X0_CG N_AI_XI2.X0_PGD 8.63152e-19
cc_301 N_BI_c_486_n N_AI_XI2.X0_PGD 0.00133285f
cc_302 N_BI_c_464_n N_AI_c_529_n 3.64122e-19
cc_303 N_BI_c_464_n N_B_c_579_n 0.00139574f
cc_304 N_BI_c_464_n N_B_c_615_n 6.02887e-19
cc_305 N_BI_c_479_n N_B_c_615_n 3.05615e-19
cc_306 N_BI_c_478_n N_B_c_583_n 0.00178808f
cc_307 N_BI_c_467_n N_B_c_583_n 0.00156529f
cc_308 N_BI_c_464_n N_B_c_620_n 4.56568e-19
cc_309 N_BI_c_486_n N_B_c_620_n 0.00266354f
cc_310 N_BI_c_487_n N_B_c_620_n 7.16621e-19
cc_311 N_BI_c_478_n N_B_c_621_n 4.56568e-19
cc_312 N_BI_c_486_n N_B_c_621_n 6.17967e-19
cc_313 N_BI_c_487_n N_B_c_621_n 0.00243716f
cc_314 N_BI_c_464_n N_B_c_581_n 0.00427216f
cc_315 N_BI_c_464_n N_B_c_603_n 3.15526e-19
cc_316 N_BI_c_467_n N_B_c_603_n 0.00129112f
cc_317 N_BI_c_506_p N_B_c_603_n 0.0034245f
cc_318 N_BI_c_464_n N_B_c_585_n 4.99817e-19
cc_319 N_BI_c_467_n N_B_c_585_n 7.12768e-19
cc_320 N_BI_c_479_n N_B_c_585_n 7.15853e-19
cc_321 N_BI_c_506_p N_B_c_645_n 0.00229162f
cc_322 N_BI_c_464_n N_B_c_586_n 0.00139788f
cc_323 N_BI_c_467_n N_B_c_586_n 8.65145e-19
cc_324 N_BI_c_464_n N_Z_c_669_n 0.00138937f
cc_325 N_BI_c_478_n N_Z_c_669_n 0.00157561f
cc_326 N_BI_c_486_n N_Z_c_669_n 8.66889e-19
cc_327 N_BI_c_467_n N_Z_c_669_n 0.00100271f
cc_328 N_BI_c_506_p N_Z_c_669_n 0.00210866f
cc_329 N_BI_c_479_n N_Z_c_669_n 9.67357e-19
cc_330 N_AI_XI2.X0_PGD N_B_c_648_n 8.79767e-19
cc_331 N_AI_c_527_n N_B_c_648_n 0.00234569f
cc_332 N_AI_c_537_n N_B_c_615_n 5.49665e-19
cc_333 N_AI_c_527_n N_B_c_615_n 4.745e-19
cc_334 N_AI_XI2.X0_PGD N_B_c_620_n 0.00133285f
cc_335 N_AI_c_566_p N_B_c_620_n 7.60534e-19
cc_336 N_AI_c_537_n N_B_c_620_n 4.46045e-19
cc_337 N_AI_c_527_n N_B_c_620_n 0.00166302f
cc_338 N_AI_c_528_n N_B_c_581_n 0.00120142f
cc_339 N_AI_c_529_n N_B_c_581_n 3.28172e-19
cc_340 N_AI_c_529_n N_B_c_602_n 2.8335e-19
cc_341 N_AI_c_537_n N_B_c_603_n 4.27113e-19
cc_342 N_AI_XI2.X0_PGD N_Z_c_669_n 3.26804e-19
cc_343 N_B_c_615_n N_Z_c_669_n 0.0013937f
cc_344 N_B_c_583_n N_Z_c_669_n 0.00139745f
cc_345 N_B_c_620_n N_Z_c_669_n 8.66889e-19
cc_346 N_B_c_621_n N_Z_c_669_n 8.66889e-19
cc_347 N_B_c_603_n N_Z_c_669_n 4.72173e-19
*
.ends
*
*
.subckt XOR3_HPNW1 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XOR3_N1
.ends
*
* File: G3_AND2_N1.pex.netlist
* Created: Wed Feb 23 10:37:48 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*






.subckt G3_AND2_N1_2 VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI7.X0 N_NET1_XI7.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_B_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW4
XI8.X0 N_NET1_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI9.X0 N_NET1_XI8.X0_D N_VSS_XI9.X0_PGD N_B_XI9.X0_CG N_VSS_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW4
XI2.X0 N_Z_XI2.X0_D N_VSS_XI2.X0_PGD N_NET1_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW4
XI1.X0 N_Z_XI2.X0_D N_VDD_XI1.X0_PGD N_NET1_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
*
x_PM_G3_AND2_N1_VSS N_VSS_XI7.X0_S N_VSS_XI8.X0_PGD N_VSS_XI8.X0_PGS
+ N_VSS_XI9.X0_PGD N_VSS_XI9.X0_PGS N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI1.X0_S N_VSS_c_13_p N_VSS_c_14_p N_VSS_c_42_p N_VSS_c_2_p N_VSS_c_49_p
+ N_VSS_c_4_p N_VSS_c_7_p N_VSS_c_23_p N_VSS_c_65_p N_VSS_c_8_p N_VSS_c_25_p
+ N_VSS_c_5_p N_VSS_c_6_p N_VSS_c_17_p N_VSS_c_10_p N_VSS_c_18_p N_VSS_c_30_p
+ N_VSS_c_68_p N_VSS_c_33_p N_VSS_c_19_p N_VSS_c_31_p VSS Vss PM_G3_AND2_N1_VSS
x_PM_G3_AND2_N1_VDD N_VDD_XI7.X0_PGD N_VDD_XI8.X0_S N_VDD_XI9.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_c_143_p N_VDD_c_128_p N_VDD_c_70_n
+ N_VDD_c_71_n N_VDD_c_75_n N_VDD_c_79_n N_VDD_c_80_n N_VDD_c_81_n N_VDD_c_116_p
+ N_VDD_c_88_n N_VDD_c_94_n N_VDD_c_100_n N_VDD_c_102_n VDD N_VDD_c_103_n
+ N_VDD_c_113_p N_VDD_c_104_n Vss PM_G3_AND2_N1_VDD
x_PM_G3_AND2_N1_A N_A_XI7.X0_CG N_A_XI8.X0_CG N_A_c_164_n N_A_c_156_n
+ N_A_c_157_n A N_A_c_167_n N_A_c_160_n Vss PM_G3_AND2_N1_A
x_PM_G3_AND2_N1_NET1 N_NET1_XI7.X0_D N_NET1_XI8.X0_D N_NET1_XI2.X0_CG
+ N_NET1_XI1.X0_CG N_NET1_c_183_n N_NET1_c_184_n N_NET1_c_185_n N_NET1_c_187_n
+ N_NET1_c_190_n N_NET1_c_193_n N_NET1_c_195_n Vss PM_G3_AND2_N1_NET1
x_PM_G3_AND2_N1_B N_B_XI7.X0_PGS N_B_XI9.X0_CG N_B_c_232_n N_B_c_234_n
+ N_B_c_239_n B N_B_c_242_n Vss PM_G3_AND2_N1_B
x_PM_G3_AND2_N1_Z N_Z_XI2.X0_D Z N_Z_c_260_n Vss PM_G3_AND2_N1_Z
cc_1 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.0016786f
cc_2 N_VSS_c_2_p N_VDD_c_70_n 0.0016786f
cc_3 N_VSS_XI7.X0_S N_VDD_c_71_n 9.73142e-19
cc_4 N_VSS_c_4_p N_VDD_c_71_n 0.0016649f
cc_5 N_VSS_c_5_p N_VDD_c_71_n 0.00583639f
cc_6 N_VSS_c_6_p N_VDD_c_71_n 0.00213268f
cc_7 N_VSS_c_7_p N_VDD_c_75_n 9.61646e-19
cc_8 N_VSS_c_8_p N_VDD_c_75_n 4.3619e-19
cc_9 N_VSS_c_5_p N_VDD_c_75_n 0.00351219f
cc_10 N_VSS_c_10_p N_VDD_c_75_n 0.00128683f
cc_11 N_VSS_c_4_p N_VDD_c_79_n 0.00221042f
cc_12 N_VSS_c_4_p N_VDD_c_80_n 7.48389e-19
cc_13 N_VSS_c_13_p N_VDD_c_81_n 0.00144388f
cc_14 N_VSS_c_14_p N_VDD_c_81_n 2.81922e-19
cc_15 N_VSS_c_7_p N_VDD_c_81_n 0.00161703f
cc_16 N_VSS_c_8_p N_VDD_c_81_n 2.03837e-19
cc_17 N_VSS_c_17_p N_VDD_c_81_n 0.00338232f
cc_18 N_VSS_c_18_p N_VDD_c_81_n 0.00635521f
cc_19 N_VSS_c_19_p N_VDD_c_81_n 7.61747e-19
cc_20 N_VSS_XI9.X0_PGS N_VDD_c_88_n 2.28184e-19
cc_21 N_VSS_XI2.X0_PGS N_VDD_c_88_n 2.56778e-19
cc_22 N_VSS_c_7_p N_VDD_c_88_n 5.65664e-19
cc_23 N_VSS_c_23_p N_VDD_c_88_n 0.00181281f
cc_24 N_VSS_c_8_p N_VDD_c_88_n 2.30125e-19
cc_25 N_VSS_c_25_p N_VDD_c_88_n 9.55109e-19
cc_26 N_VSS_c_2_p N_VDD_c_94_n 4.8598e-19
cc_27 N_VSS_c_23_p N_VDD_c_94_n 0.00161703f
cc_28 N_VSS_c_25_p N_VDD_c_94_n 2.03837e-19
cc_29 N_VSS_c_18_p N_VDD_c_94_n 0.00145178f
cc_30 N_VSS_c_30_p N_VDD_c_94_n 0.00590089f
cc_31 N_VSS_c_31_p N_VDD_c_94_n 7.74609e-19
cc_32 N_VSS_c_23_p N_VDD_c_100_n 8.94411e-19
cc_33 N_VSS_c_33_p N_VDD_c_100_n 3.85245e-19
cc_34 N_VSS_c_5_p N_VDD_c_102_n 0.00104993f
cc_35 N_VSS_c_18_p N_VDD_c_103_n 0.00119068f
cc_36 N_VSS_c_23_p N_VDD_c_104_n 3.48267e-19
cc_37 N_VSS_c_25_p N_VDD_c_104_n 8.0279e-19
cc_38 N_VSS_c_8_p N_A_c_156_n 0.00234241f
cc_39 N_VSS_c_7_p N_A_c_157_n 8.12473e-19
cc_40 N_VSS_c_8_p N_A_c_157_n 5.42695e-19
cc_41 N_VSS_c_5_p N_A_c_157_n 6.55807e-19
cc_42 N_VSS_c_42_p N_A_c_160_n 7.84334e-19
cc_43 N_VSS_c_7_p N_A_c_160_n 4.56568e-19
cc_44 N_VSS_c_8_p N_A_c_160_n 0.00184767f
cc_45 N_VSS_XI7.X0_S N_NET1_XI7.X0_D 3.43419e-19
cc_46 N_VSS_c_4_p N_NET1_XI7.X0_D 3.48267e-19
cc_47 N_VSS_c_25_p N_NET1_c_183_n 0.00413078f
cc_48 N_VSS_XI2.X0_PGD N_NET1_c_184_n 4.20799e-19
cc_49 N_VSS_c_49_p N_NET1_c_185_n 9.28737e-19
cc_50 N_VSS_c_25_p N_NET1_c_185_n 2.03369e-19
cc_51 N_VSS_XI7.X0_S N_NET1_c_187_n 3.48267e-19
cc_52 N_VSS_c_4_p N_NET1_c_187_n 8.46599e-19
cc_53 N_VSS_c_5_p N_NET1_c_187_n 2.07501e-19
cc_54 N_VSS_c_23_p N_NET1_c_190_n 0.00125323f
cc_55 N_VSS_c_25_p N_NET1_c_190_n 4.64764e-19
cc_56 N_VSS_c_5_p N_NET1_c_190_n 3.39684e-19
cc_57 N_VSS_c_23_p N_NET1_c_193_n 4.56568e-19
cc_58 N_VSS_c_25_p N_NET1_c_193_n 6.1245e-19
cc_59 N_VSS_c_5_p N_NET1_c_195_n 2.06399e-19
cc_60 N_VSS_c_18_p N_NET1_c_195_n 0.00149275f
cc_61 N_VSS_XI8.X0_PGD N_B_c_232_n 6.72196e-19
cc_62 N_VSS_XI9.X0_PGD N_B_c_232_n 6.72196e-19
cc_63 N_VSS_XI8.X0_PGS N_B_c_234_n 7.85613e-19
cc_64 N_VSS_XI1.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_65 N_VSS_c_65_p N_Z_XI2.X0_D 3.48267e-19
cc_66 N_VSS_c_65_p N_Z_c_260_n 5.37696e-19
cc_67 N_VSS_c_30_p N_Z_c_260_n 2.64173e-19
cc_68 N_VSS_c_68_p N_Z_c_260_n 2.7826e-19
cc_69 N_VDD_XI7.X0_PGD N_A_XI7.X0_CG 4.88425e-19
cc_70 N_VDD_c_79_n N_A_c_164_n 3.72495e-19
cc_71 N_VDD_c_71_n N_A_c_157_n 0.00273528f
cc_72 N_VDD_c_79_n N_A_c_157_n 7.03725e-19
cc_73 N_VDD_XI7.X0_PGD N_A_c_167_n 2.88617e-19
cc_74 N_VDD_c_71_n N_A_c_167_n 3.68786e-19
cc_75 N_VDD_c_79_n N_A_c_167_n 4.3265e-19
cc_76 N_VDD_c_113_p N_A_c_167_n 7.96439e-19
cc_77 N_VDD_c_71_n N_A_c_160_n 5.09899e-19
cc_78 N_VDD_c_79_n N_NET1_XI7.X0_D 9.18655e-19
cc_79 N_VDD_c_116_p N_NET1_XI7.X0_D 8.835e-19
cc_80 N_VDD_c_113_p N_NET1_XI7.X0_D 0.00132057f
cc_81 N_VDD_XI8.X0_S N_NET1_XI8.X0_D 3.43419e-19
cc_82 N_VDD_XI9.X0_S N_NET1_XI8.X0_D 3.43419e-19
cc_83 N_VDD_c_80_n N_NET1_XI8.X0_D 3.74351e-19
cc_84 N_VDD_c_81_n N_NET1_XI8.X0_D 3.7884e-19
cc_85 N_VDD_c_88_n N_NET1_XI8.X0_D 3.48267e-19
cc_86 N_VDD_c_104_n N_NET1_XI1.X0_CG 8.03148e-19
cc_87 N_VDD_XI1.X0_PGD N_NET1_c_184_n 4.25379e-19
cc_88 N_VDD_XI7.X0_PGD N_NET1_c_187_n 2.94751e-19
cc_89 N_VDD_XI8.X0_S N_NET1_c_187_n 3.48267e-19
cc_90 N_VDD_XI9.X0_S N_NET1_c_187_n 3.48267e-19
cc_91 N_VDD_c_128_p N_NET1_c_187_n 5.10453e-19
cc_92 N_VDD_c_71_n N_NET1_c_187_n 6.49505e-19
cc_93 N_VDD_c_79_n N_NET1_c_187_n 0.00151981f
cc_94 N_VDD_c_80_n N_NET1_c_187_n 8.1398e-19
cc_95 N_VDD_c_81_n N_NET1_c_187_n 5.36364e-19
cc_96 N_VDD_c_116_p N_NET1_c_187_n 0.00366419f
cc_97 N_VDD_c_88_n N_NET1_c_187_n 7.99681e-19
cc_98 N_VDD_c_113_p N_NET1_c_187_n 8.835e-19
cc_99 N_VDD_c_79_n N_NET1_c_195_n 3.89533e-19
cc_100 N_VDD_c_81_n N_NET1_c_195_n 3.69547e-19
cc_101 N_VDD_c_116_p N_NET1_c_195_n 4.83374e-19
cc_102 N_VDD_c_88_n N_NET1_c_195_n 4.34102e-19
cc_103 N_VDD_XI7.X0_PGD N_B_XI7.X0_PGS 0.00320719f
cc_104 N_VDD_c_71_n N_B_XI7.X0_PGS 6.17633e-19
cc_105 N_VDD_c_79_n N_B_XI7.X0_PGS 2.2956e-19
cc_106 N_VDD_c_143_p N_B_c_232_n 0.00973324f
cc_107 N_VDD_c_81_n N_B_c_239_n 4.48125e-19
cc_108 N_VDD_c_116_p N_B_c_239_n 4.13122e-19
cc_109 N_VDD_c_113_p N_B_c_239_n 0.00150022f
cc_110 N_VDD_c_81_n N_B_c_242_n 2.66883e-19
cc_111 N_VDD_c_116_p N_B_c_242_n 3.55986e-19
cc_112 N_VDD_c_113_p N_B_c_242_n 3.81676e-19
cc_113 N_VDD_XI9.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_114 N_VDD_c_88_n N_Z_XI2.X0_D 3.48267e-19
cc_115 N_VDD_c_94_n N_Z_XI2.X0_D 3.7884e-19
cc_116 N_VDD_XI9.X0_S N_Z_c_260_n 3.48267e-19
cc_117 N_VDD_c_88_n N_Z_c_260_n 7.06424e-19
cc_118 N_VDD_c_94_n N_Z_c_260_n 5.12447e-19
cc_119 N_A_c_157_n N_NET1_c_187_n 0.00751692f
cc_120 N_A_c_167_n N_NET1_c_187_n 9.57699e-19
cc_121 N_A_c_160_n N_NET1_c_187_n 9.18163e-19
cc_122 N_A_XI7.X0_CG N_B_XI7.X0_PGS 4.5346e-19
cc_123 N_A_c_167_n N_B_XI7.X0_PGS 5.70584e-19
cc_124 N_A_c_157_n N_B_c_232_n 2.1473e-19
cc_125 N_A_c_167_n N_B_c_232_n 0.0014179f
cc_126 N_A_c_160_n N_B_c_232_n 0.00112482f
cc_127 N_A_c_160_n N_B_c_239_n 9.27569e-19
cc_128 N_NET1_c_187_n N_B_c_232_n 7.63501e-19
cc_129 N_NET1_c_187_n N_B_c_239_n 9.91045e-19
cc_130 N_NET1_c_190_n N_B_c_239_n 3.63713e-19
cc_131 N_NET1_c_193_n N_B_c_239_n 0.00197331f
cc_132 N_NET1_c_187_n N_B_c_242_n 0.00142922f
cc_133 N_NET1_c_190_n N_B_c_242_n 3.90886e-19
cc_134 N_NET1_c_193_n N_B_c_242_n 3.48267e-19
*
.ends
*
*
.subckt AND2_HPNW4 A B Y VDD VSS
xgate (VSS VDD A B Y) G3_AND2_N1_2
.ends
*
* File: G2_AOI21_N1.pex.netlist
* Created: Mon Apr 11 11:24:15 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*






.subckt G2_AOI21_N1_2 VSS VDD B C Z A
*
* A	A
* Z	Z
* C	C
* B	B
* VDD	VDD
* VSS	VSS
XI1.X0 N_Z_XI1.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_B_XI1.X0_PGS N_VSS_XI1.X0_S
+ TIGFET_HPNW4
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_C_XI6.X0_PGS N_VDD_XI6.X0_S
+ TIGFET_HPNW4
XI5.X0 N_Z_XI1.X0_D N_VDD_XI5.X0_PGD N_C_XI5.X0_CG N_VDD_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW4
XI7.X0 N_Z_XI6.X0_D N_VSS_XI7.X0_PGD N_A_XI7.X0_CG N_C_XI7.X0_PGS N_VDD_XI7.X0_S
+ TIGFET_HPNW4
*
x_PM_G2_AOI21_N1_VSS N_VSS_XI1.X0_S N_VSS_XI6.X0_PGD N_VSS_XI5.X0_S
+ N_VSS_XI7.X0_PGD N_VSS_c_3_p N_VSS_c_46_p N_VSS_c_2_p N_VSS_c_4_p N_VSS_c_8_p
+ N_VSS_c_20_p N_VSS_c_23_p N_VSS_c_9_p N_VSS_c_1_p N_VSS_c_5_p N_VSS_c_6_p
+ N_VSS_c_13_p N_VSS_c_10_p N_VSS_c_16_p N_VSS_c_17_p VSS N_VSS_c_18_p Vss
+ PM_G2_AOI21_N1_VSS
x_PM_G2_AOI21_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI6.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI5.X0_PGS N_VDD_XI7.X0_S N_VDD_c_89_p N_VDD_c_54_n N_VDD_c_55_n
+ N_VDD_c_56_n N_VDD_c_77_p N_VDD_c_60_n N_VDD_c_64_n N_VDD_c_65_n N_VDD_c_67_n
+ N_VDD_c_72_n VDD N_VDD_c_75_n N_VDD_c_78_p Vss PM_G2_AOI21_N1_VDD
x_PM_G2_AOI21_N1_B N_B_XI1.X0_PGS N_B_XI6.X0_CG N_B_c_122_p B N_B_c_119_n Vss
+ PM_G2_AOI21_N1_B
x_PM_G2_AOI21_N1_C N_C_XI6.X0_PGS N_C_XI5.X0_CG N_C_XI7.X0_PGS N_C_c_143_n
+ N_C_c_146_n N_C_c_147_n N_C_c_134_n C N_C_c_136_n C N_C_c_137_n N_C_c_140_n
+ Vss PM_G2_AOI21_N1_C
x_PM_G2_AOI21_N1_Z N_Z_XI1.X0_D N_Z_XI6.X0_D N_Z_c_182_n Z Vss PM_G2_AOI21_N1_Z
x_PM_G2_AOI21_N1_A N_A_XI1.X0_CG N_A_XI7.X0_CG N_A_c_208_n N_A_c_225_n
+ N_A_c_226_n N_A_c_209_n N_A_c_227_n N_A_c_211_n N_A_c_212_n A N_A_c_216_n Vss
+ PM_G2_AOI21_N1_A
cc_1 N_VSS_c_1_p N_VDD_c_54_n 4.93612e-19
cc_2 N_VSS_c_2_p N_VDD_c_55_n 9.30121e-19
cc_3 N_VSS_c_3_p N_VDD_c_56_n 0.0011834f
cc_4 N_VSS_c_4_p N_VDD_c_56_n 0.00161703f
cc_5 N_VSS_c_5_p N_VDD_c_56_n 0.00445263f
cc_6 N_VSS_c_6_p N_VDD_c_56_n 0.00169823f
cc_7 N_VSS_XI5.X0_S N_VDD_c_60_n 3.83684e-19
cc_8 N_VSS_c_8_p N_VDD_c_60_n 4.79306e-19
cc_9 N_VSS_c_9_p N_VDD_c_60_n 0.0035571f
cc_10 N_VSS_c_10_p N_VDD_c_60_n 0.00109026f
cc_11 N_VSS_c_9_p N_VDD_c_64_n 0.00162315f
cc_12 N_VSS_c_8_p N_VDD_c_65_n 2.13058e-19
cc_13 N_VSS_c_13_p N_VDD_c_65_n 5.33968e-19
cc_14 N_VSS_XI5.X0_S N_VDD_c_67_n 9.5668e-19
cc_15 N_VSS_c_8_p N_VDD_c_67_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_67_n 0.00300233f
cc_17 N_VSS_c_17_p N_VDD_c_67_n 0.00605714f
cc_18 N_VSS_c_18_p N_VDD_c_67_n 8.91588e-19
cc_19 N_VSS_c_4_p N_VDD_c_72_n 4.42697e-19
cc_20 N_VSS_c_20_p N_VDD_c_72_n 3.70842e-19
cc_21 N_VSS_c_17_p N_VDD_c_72_n 0.00278561f
cc_22 N_VSS_c_17_p N_VDD_c_75_n 9.45256e-19
cc_23 N_VSS_c_23_p B 3.22996e-19
cc_24 N_VSS_c_9_p B 3.31649e-19
cc_25 N_VSS_XI6.X0_PGD N_C_XI6.X0_PGS 0.00161425f
cc_26 N_VSS_c_4_p N_C_c_134_n 5.88052e-19
cc_27 N_VSS_c_17_p N_C_c_134_n 0.00138265f
cc_28 N_VSS_c_17_p N_C_c_136_n 3.65158e-19
cc_29 N_VSS_XI6.X0_PGD N_C_c_137_n 3.23173e-19
cc_30 N_VSS_c_4_p N_C_c_137_n 3.44698e-19
cc_31 N_VSS_c_20_p N_C_c_137_n 3.34921e-19
cc_32 N_VSS_c_9_p N_C_c_140_n 0.00303126f
cc_33 N_VSS_c_17_p N_C_c_140_n 3.90377e-19
cc_34 N_VSS_XI1.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_35 N_VSS_XI5.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_XI1.X0_D 3.48267e-19
cc_37 N_VSS_c_8_p N_Z_XI1.X0_D 3.48267e-19
cc_38 N_VSS_XI1.X0_S N_Z_c_182_n 3.48267e-19
cc_39 N_VSS_XI5.X0_S N_Z_c_182_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_182_n 5.69026e-19
cc_41 N_VSS_c_8_p N_Z_c_182_n 5.69026e-19
cc_42 N_VSS_c_9_p N_Z_c_182_n 4.18012e-19
cc_43 N_VSS_c_17_p N_Z_c_182_n 5.20852e-19
cc_44 N_VSS_XI6.X0_PGD N_A_c_208_n 7.38139e-19
cc_45 N_VSS_XI7.X0_PGD N_A_c_209_n 0.00160007f
cc_46 N_VSS_c_46_p N_A_c_209_n 3.07681e-19
cc_47 N_VSS_c_20_p N_A_c_211_n 0.00255152f
cc_48 N_VSS_c_46_p N_A_c_212_n 8.89952e-19
cc_49 N_VSS_c_20_p N_A_c_212_n 2.75949e-19
cc_50 N_VSS_c_4_p A 5.37794e-19
cc_51 N_VSS_c_20_p A 4.56568e-19
cc_52 N_VSS_c_4_p N_A_c_216_n 4.56568e-19
cc_53 N_VSS_c_20_p N_A_c_216_n 6.1245e-19
cc_54 N_VDD_XI1.X0_PGD N_B_XI1.X0_PGS 0.0015605f
cc_55 N_VDD_c_77_p B 5.21626e-19
cc_56 N_VDD_c_78_p B 3.48267e-19
cc_57 N_VDD_XI1.X0_PGD N_B_c_119_n 3.73456e-19
cc_58 N_VDD_c_77_p N_B_c_119_n 4.2695e-19
cc_59 N_VDD_c_78_p N_B_c_119_n 5.71625e-19
cc_60 N_VDD_c_78_p N_C_XI5.X0_CG 0.00117555f
cc_61 N_VDD_c_77_p N_C_c_143_n 4.85469e-19
cc_62 N_VDD_c_67_n N_C_c_143_n 5.82627e-19
cc_63 N_VDD_c_78_p N_C_c_143_n 0.00182135f
cc_64 N_VDD_c_56_n N_C_c_146_n 3.54083e-19
cc_65 N_VDD_XI5.X0_PGS N_C_c_147_n 7.91098e-19
cc_66 N_VDD_c_67_n N_C_c_147_n 4.33233e-19
cc_67 N_VDD_c_89_p N_C_c_134_n 3.48763e-19
cc_68 N_VDD_c_55_n N_C_c_134_n 3.25844e-19
cc_69 N_VDD_c_56_n N_C_c_134_n 0.00156477f
cc_70 N_VDD_c_56_n N_C_c_136_n 7.40864e-19
cc_71 N_VDD_c_77_p N_C_c_136_n 5.82566e-19
cc_72 N_VDD_c_67_n N_C_c_136_n 4.90875e-19
cc_73 N_VDD_c_78_p N_C_c_136_n 4.56568e-19
cc_74 N_VDD_c_89_p N_C_c_137_n 4.55865e-19
cc_75 N_VDD_c_56_n N_C_c_137_n 2.55177e-19
cc_76 N_VDD_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_77 N_VDD_XI7.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_78 N_VDD_c_55_n N_Z_XI6.X0_D 3.72199e-19
cc_79 N_VDD_c_56_n N_Z_XI6.X0_D 3.7884e-19
cc_80 N_VDD_c_65_n N_Z_XI6.X0_D 3.72199e-19
cc_81 N_VDD_XI6.X0_S N_Z_c_182_n 3.48267e-19
cc_82 N_VDD_XI7.X0_S N_Z_c_182_n 3.48267e-19
cc_83 N_VDD_c_55_n N_Z_c_182_n 5.68773e-19
cc_84 N_VDD_c_56_n N_Z_c_182_n 6.9352e-19
cc_85 N_VDD_c_65_n N_Z_c_182_n 7.77875e-19
cc_86 N_VDD_c_67_n N_Z_c_182_n 9.95668e-19
cc_87 N_VDD_XI1.X0_PGD N_A_c_208_n 6.1925e-19
cc_88 N_VDD_XI5.X0_PGD N_A_c_209_n 3.67852e-19
cc_89 N_VDD_c_67_n A 3.35548e-19
cc_90 N_VDD_c_56_n N_A_c_216_n 2.29043e-19
cc_91 N_VDD_c_67_n N_A_c_216_n 3.66936e-19
cc_92 N_B_c_122_p N_C_XI6.X0_PGS 0.00189436f
cc_93 N_B_XI1.X0_PGS N_C_XI5.X0_CG 2.46172e-19
cc_94 N_B_c_122_p N_C_XI7.X0_PGS 4.95875e-19
cc_95 N_B_c_122_p N_C_c_146_n 3.12087e-19
cc_96 N_B_XI1.X0_PGS N_Z_c_182_n 2.61881e-19
cc_97 N_B_XI1.X0_PGS N_A_XI1.X0_CG 0.00900711f
cc_98 N_B_c_119_n N_A_XI1.X0_CG 0.00150571f
cc_99 N_B_c_122_p N_A_c_225_n 0.00163406f
cc_100 N_B_XI1.X0_PGS N_A_c_226_n 6.07734e-19
cc_101 N_B_c_122_p N_A_c_227_n 0.00136506f
cc_102 N_B_c_122_p N_A_c_216_n 2.87722e-19
cc_103 N_C_c_143_n N_Z_c_182_n 9.29334e-19
cc_104 N_C_c_134_n N_Z_c_182_n 0.00223036f
cc_105 N_C_c_136_n N_Z_c_182_n 0.00299789f
cc_106 N_C_c_140_n N_Z_c_182_n 2.70867e-19
cc_107 N_C_XI5.X0_CG N_A_XI1.X0_CG 5.49495e-19
cc_108 N_C_c_143_n N_A_XI1.X0_CG 5.65259e-19
cc_109 N_C_XI7.X0_PGS N_A_c_208_n 8.10159e-19
cc_110 N_C_c_147_n N_A_c_208_n 0.00121323f
cc_111 N_C_XI7.X0_PGS N_A_c_211_n 5.00154e-19
cc_112 N_C_c_143_n N_A_c_212_n 9.55393e-19
cc_113 N_C_c_143_n A 4.56568e-19
cc_114 N_C_c_136_n A 6.2998e-19
cc_115 N_C_XI7.X0_PGS N_A_c_216_n 0.00570455f
cc_116 N_C_c_143_n N_A_c_216_n 8.77002e-19
cc_117 N_C_c_147_n N_A_c_216_n 0.00119367f
cc_118 N_C_c_136_n N_A_c_216_n 4.56568e-19
cc_119 N_Z_c_182_n N_A_XI1.X0_CG 5.75111e-19
cc_120 N_Z_c_182_n N_A_c_208_n 4.34888e-19
cc_121 N_Z_c_182_n A 0.0015179f
cc_122 N_Z_c_182_n N_A_c_216_n 8.99071e-19
*
.ends
*
*
.subckt AOI21_HPNW4 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 B0 Y A0) G2_AOI21_N1_2
.ends
*
* File: G2_BUF1_N1.pex.netlist
* Created: Wed Mar  2 15:26:00 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*





.subckt G2_BUF1_N1_2 VDD VSS A Z
*
* Z	Z
* A	A
* VSS	VSS
* VDD	VDD
XI3.X0 N_Z_XI3.X0_D N_VSS_XI3.X0_PGD N_NET17_XI3.X0_CG N_VSS_XI3.X0_PGD
+ N_VDD_XI3.X0_S TIGFET_HPNW4
XI2.X0 N_NET17_XI2.X0_D N_VSS_XI2.X0_PGD N_A_XI2.X0_CG N_VSS_XI2.X0_PGD
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI0.X0 N_Z_XI3.X0_D N_VDD_XI0.X0_PGD N_NET17_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW4
XI1.X0 N_NET17_XI2.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW4
*
x_PM_G2_BUF1_N1_VDD N_VDD_XI3.X0_S N_VDD_XI2.X0_S N_VDD_XI0.X0_PGD
+ N_VDD_XI1.X0_PGD N_VDD_c_3_p N_VDD_c_6_p N_VDD_c_9_p VDD N_VDD_c_13_p
+ N_VDD_c_4_p N_VDD_c_38_p N_VDD_c_43_p N_VDD_c_7_p N_VDD_c_11_p N_VDD_c_15_p
+ N_VDD_c_12_p N_VDD_c_16_p Vss PM_G2_BUF1_N1_VDD
x_PM_G2_BUF1_N1_VSS N_VSS_XI3.X0_PGD N_VSS_XI2.X0_PGD N_VSS_XI0.X0_S
+ N_VSS_XI1.X0_S N_VSS_c_61_n N_VSS_c_63_n N_VSS_c_64_n N_VSS_c_66_n
+ N_VSS_c_67_n N_VSS_c_71_n N_VSS_c_101_p N_VSS_c_110_p N_VSS_c_75_n
+ N_VSS_c_79_n N_VSS_c_83_n N_VSS_c_84_n N_VSS_c_85_n N_VSS_c_86_n N_VSS_c_104_p
+ N_VSS_c_112_p N_VSS_c_87_n VSS N_VSS_c_88_n Vss PM_G2_BUF1_N1_VSS
x_PM_G2_BUF1_N1_A N_A_XI2.X0_CG N_A_XI1.X0_CG N_A_c_124_n N_A_c_120_n A
+ N_A_c_122_n N_A_c_123_n Vss PM_G2_BUF1_N1_A
x_PM_G2_BUF1_N1_Z N_Z_XI3.X0_D Z Vss PM_G2_BUF1_N1_Z
x_PM_G2_BUF1_N1_NET17 N_NET17_XI3.X0_CG N_NET17_XI2.X0_D N_NET17_XI0.X0_CG
+ N_NET17_c_155_n N_NET17_c_157_n N_NET17_c_160_n N_NET17_c_164_n
+ N_NET17_c_168_n Vss PM_G2_BUF1_N1_NET17
cc_1 N_VDD_XI0.X0_PGD N_VSS_XI3.X0_PGD 0.00173038f
cc_2 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00173038f
cc_3 N_VDD_c_3_p N_VSS_c_61_n 0.00173038f
cc_4 N_VDD_c_4_p N_VSS_c_61_n 2.91357e-19
cc_5 N_VDD_c_4_p N_VSS_c_63_n 3.24852e-19
cc_6 N_VDD_c_6_p N_VSS_c_64_n 0.00173038f
cc_7 N_VDD_c_7_p N_VSS_c_64_n 2.91357e-19
cc_8 N_VDD_c_7_p N_VSS_c_66_n 3.24852e-19
cc_9 N_VDD_c_9_p N_VSS_c_67_n 8.69498e-19
cc_10 N_VDD_c_4_p N_VSS_c_67_n 0.00141228f
cc_11 N_VDD_c_11_p N_VSS_c_67_n 0.00106872f
cc_12 N_VDD_c_12_p N_VSS_c_67_n 3.48267e-19
cc_13 N_VDD_c_13_p N_VSS_c_71_n 8.69498e-19
cc_14 N_VDD_c_7_p N_VSS_c_71_n 0.00141228f
cc_15 N_VDD_c_15_p N_VSS_c_71_n 0.00106872f
cc_16 N_VDD_c_16_p N_VSS_c_71_n 3.48267e-19
cc_17 N_VDD_c_9_p N_VSS_c_75_n 3.66936e-19
cc_18 N_VDD_c_4_p N_VSS_c_75_n 0.00112249f
cc_19 N_VDD_c_11_p N_VSS_c_75_n 3.99794e-19
cc_20 N_VDD_c_12_p N_VSS_c_75_n 8.09245e-19
cc_21 N_VDD_c_13_p N_VSS_c_79_n 3.66936e-19
cc_22 N_VDD_c_7_p N_VSS_c_79_n 0.00112249f
cc_23 N_VDD_c_15_p N_VSS_c_79_n 3.99794e-19
cc_24 N_VDD_c_16_p N_VSS_c_79_n 8.09245e-19
cc_25 N_VDD_c_4_p N_VSS_c_83_n 0.00554293f
cc_26 N_VDD_c_4_p N_VSS_c_84_n 0.0017359f
cc_27 N_VDD_c_7_p N_VSS_c_85_n 0.00562924f
cc_28 N_VDD_c_7_p N_VSS_c_86_n 0.0017359f
cc_29 N_VDD_c_11_p N_VSS_c_87_n 3.85245e-19
cc_30 N_VDD_c_15_p N_VSS_c_88_n 3.85245e-19
cc_31 N_VDD_c_16_p N_A_XI1.X0_CG 0.00254294f
cc_32 N_VDD_XI0.X0_PGD N_A_c_120_n 4.08785e-19
cc_33 N_VDD_XI1.X0_PGD N_A_c_120_n 4.04053e-19
cc_34 VDD N_A_c_122_n 5.94555e-19
cc_35 VDD N_A_c_123_n 4.56718e-19
cc_36 N_VDD_XI3.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_37 N_VDD_c_4_p N_Z_XI3.X0_D 3.7884e-19
cc_38 N_VDD_c_38_p N_Z_XI3.X0_D 3.72199e-19
cc_39 N_VDD_XI3.X0_S Z 3.48267e-19
cc_40 N_VDD_c_4_p Z 5.12447e-19
cc_41 N_VDD_c_38_p Z 7.4527e-19
cc_42 N_VDD_XI2.X0_S N_NET17_XI2.X0_D 3.43419e-19
cc_43 N_VDD_c_43_p N_NET17_XI2.X0_D 3.72199e-19
cc_44 N_VDD_c_12_p N_NET17_XI0.X0_CG 0.0023817f
cc_45 N_VDD_XI0.X0_PGD N_NET17_c_155_n 4.04053e-19
cc_46 N_VDD_XI1.X0_PGD N_NET17_c_155_n 4.08785e-19
cc_47 N_VDD_XI2.X0_S N_NET17_c_157_n 3.48267e-19
cc_48 N_VDD_c_43_p N_NET17_c_157_n 8.0086e-19
cc_49 N_VDD_c_7_p N_NET17_c_157_n 5.01863e-19
cc_50 N_VDD_c_11_p N_NET17_c_160_n 6.85072e-19
cc_51 N_VDD_c_15_p N_NET17_c_160_n 3.98507e-19
cc_52 N_VDD_c_12_p N_NET17_c_160_n 4.99367e-19
cc_53 N_VDD_c_16_p N_NET17_c_160_n 3.0441e-19
cc_54 N_VDD_c_11_p N_NET17_c_164_n 4.85469e-19
cc_55 N_VDD_c_15_p N_NET17_c_164_n 3.00204e-19
cc_56 N_VDD_c_12_p N_NET17_c_164_n 0.0014909f
cc_57 N_VDD_c_16_p N_NET17_c_164_n 6.61247e-19
cc_58 VDD N_NET17_c_168_n 3.1911e-19
cc_59 N_VSS_c_79_n N_A_c_124_n 0.0023454f
cc_60 N_VSS_XI3.X0_PGD N_A_c_120_n 4.07282e-19
cc_61 N_VSS_XI2.X0_PGD N_A_c_120_n 3.99472e-19
cc_62 N_VSS_c_67_n N_A_c_122_n 2.85158e-19
cc_63 N_VSS_c_71_n N_A_c_122_n 5.53028e-19
cc_64 N_VSS_c_75_n N_A_c_122_n 3.0441e-19
cc_65 N_VSS_c_79_n N_A_c_122_n 4.99367e-19
cc_66 N_VSS_c_67_n N_A_c_123_n 2.82333e-19
cc_67 N_VSS_c_71_n N_A_c_123_n 4.56568e-19
cc_68 N_VSS_c_75_n N_A_c_123_n 6.61247e-19
cc_69 N_VSS_c_79_n N_A_c_123_n 0.0014909f
cc_70 N_VSS_XI0.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_71 N_VSS_c_101_p N_Z_XI3.X0_D 3.48267e-19
cc_72 N_VSS_XI0.X0_S Z 3.48267e-19
cc_73 N_VSS_c_101_p Z 4.99861e-19
cc_74 N_VSS_c_104_p Z 2.7826e-19
cc_75 N_VSS_c_75_n N_NET17_XI3.X0_CG 0.00250664f
cc_76 N_VSS_XI1.X0_S N_NET17_XI2.X0_D 3.43419e-19
cc_77 N_VSS_XI3.X0_PGD N_NET17_c_155_n 3.99472e-19
cc_78 N_VSS_XI2.X0_PGD N_NET17_c_155_n 4.07282e-19
cc_79 N_VSS_XI1.X0_S N_NET17_c_157_n 3.48267e-19
cc_80 N_VSS_c_110_p N_NET17_c_157_n 4.8288e-19
cc_81 N_VSS_c_85_n N_NET17_c_157_n 5.36354e-19
cc_82 N_VSS_c_112_p N_NET17_c_157_n 5.49885e-19
cc_83 VSS N_NET17_c_157_n 6.44069e-19
cc_84 N_VSS_c_83_n N_NET17_c_160_n 3.16821e-19
cc_85 N_VSS_c_85_n N_NET17_c_160_n 2.03753e-19
cc_86 VSS N_NET17_c_160_n 8.09756e-19
cc_87 N_VSS_c_83_n N_NET17_c_168_n 0.00101305f
cc_88 N_VSS_c_85_n N_NET17_c_168_n 5.70583e-19
cc_89 N_A_c_120_n N_NET17_c_155_n 0.00954069f
cc_90 N_A_c_122_n N_NET17_c_157_n 8.44937e-19
cc_91 N_Z_XI3.X0_D N_NET17_XI2.X0_D 2.56268e-19
cc_92 Z N_NET17_XI2.X0_D 3.17139e-19
cc_93 N_Z_XI3.X0_D N_NET17_c_157_n 3.17139e-19
cc_94 Z N_NET17_c_157_n 3.16516e-19
*
.ends
*
*
.subckt BUF1_HPNW4 A Y VDD VSS
xgate (VDD VSS A Y) G2_BUF1_N1_2
.ends
*
* File: G3_DFFQ1_N1.pex.netlist
* Created: Tue Apr  5 22:58:19 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*







.subckt G3_DFFQ1_N1_2 VSS CK VDD D Q
*
* Q	Q
* D	D
* VDD	VDD
* CK	CK
* VSS	VSS
XI1.X0 N_CKN_XI1.X0_D N_VDD_XI1.X0_PGD N_CK_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI2.X0 N_CKN_XI1.X0_D N_VSS_XI2.X0_PGD N_CK_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI5.X0 N_X_XI5.X0_D N_VSS_XI5.X0_PGD N_D_XI5.X0_CG N_CK_XI5.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI3.X0 N_Q_XI3.X0_D N_VDD_XI3.X0_PGD N_X_XI3.X0_CG N_CK_XI3.X0_PGS
+ N_VSS_XI3.X0_S TIGFET_HPNW4
XI4.X0 N_X_XI5.X0_D N_VDD_XI4.X0_PGD N_D_XI4.X0_CG N_CKN_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW4
XI0.X0 N_Q_XI3.X0_D N_VSS_XI0.X0_PGD N_X_XI0.X0_CG N_CKN_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW4
*
x_PM_G3_DFFQ1_N1_VSS N_VSS_XI1.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI5.X0_PGD N_VSS_XI3.X0_S N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_11_p
+ N_VSS_c_89_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_15_p N_VSS_c_3_p N_VSS_c_32_p
+ N_VSS_c_23_p N_VSS_c_33_p N_VSS_c_45_p N_VSS_c_20_p N_VSS_c_4_p N_VSS_c_34_p
+ N_VSS_c_16_p N_VSS_c_7_p N_VSS_c_22_p N_VSS_c_17_p N_VSS_c_85_p VSS
+ N_VSS_c_38_p N_VSS_c_29_p N_VSS_c_39_p N_VSS_c_48_p N_VSS_c_51_p N_VSS_c_52_p
+ N_VSS_c_30_p N_VSS_c_40_p N_VSS_c_53_p Vss PM_G3_DFFQ1_N1_VSS
x_PM_G3_DFFQ1_N1_CK N_CK_XI1.X0_CG N_CK_XI2.X0_CG N_CK_XI5.X0_PGS
+ N_CK_XI3.X0_PGS N_CK_c_122_n N_CK_c_123_n CK N_CK_c_129_p Vss
+ PM_G3_DFFQ1_N1_CK
x_PM_G3_DFFQ1_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI2.X0_S
+ N_VDD_XI3.X0_PGD N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_152_n N_VDD_c_250_p
+ N_VDD_c_153_n N_VDD_c_154_n N_VDD_c_155_n N_VDD_c_159_n N_VDD_c_163_n
+ N_VDD_c_164_n N_VDD_c_166_n N_VDD_c_172_n N_VDD_c_176_n N_VDD_c_182_n
+ N_VDD_c_183_n N_VDD_c_185_n N_VDD_c_188_n N_VDD_c_190_n N_VDD_c_195_n
+ N_VDD_c_199_n N_VDD_c_201_n N_VDD_c_203_n N_VDD_c_204_n N_VDD_c_205_n VDD
+ N_VDD_c_206_n N_VDD_c_208_n N_VDD_c_211_n Vss PM_G3_DFFQ1_N1_VDD
x_PM_G3_DFFQ1_N1_CKN N_CKN_XI1.X0_D N_CKN_XI4.X0_PGS N_CKN_XI0.X0_PGS
+ N_CKN_c_283_n N_CKN_c_268_n N_CKN_c_272_n N_CKN_c_274_n Vss PM_G3_DFFQ1_N1_CKN
x_PM_G3_DFFQ1_N1_D N_D_XI5.X0_CG N_D_XI4.X0_CG N_D_c_305_n N_D_c_306_n D
+ N_D_c_308_n N_D_c_312_n Vss PM_G3_DFFQ1_N1_D
x_PM_G3_DFFQ1_N1_X N_X_XI5.X0_D N_X_XI3.X0_CG N_X_XI0.X0_CG N_X_c_346_n
+ N_X_c_334_n N_X_c_354_n N_X_c_336_n N_X_c_337_n N_X_c_341_n N_X_c_343_n Vss
+ PM_G3_DFFQ1_N1_X
x_PM_G3_DFFQ1_N1_Q N_Q_XI3.X0_D Q Vss PM_G3_DFFQ1_N1_Q
cc_1 N_VSS_XI2.X0_PGS N_CK_XI5.X0_PGS 0.0029499f
cc_2 N_VSS_XI5.X0_PGD N_CK_XI5.X0_PGS 0.00158255f
cc_3 N_VSS_c_3_p N_CK_XI5.X0_PGS 8.20198e-19
cc_4 N_VSS_c_4_p N_CK_XI5.X0_PGS 4.62582e-19
cc_5 N_VSS_XI2.X0_PGD N_CK_c_122_n 4.16623e-19
cc_6 N_VSS_XI2.X0_PGS N_CK_c_123_n 4.26524e-19
cc_7 N_VSS_c_7_p CK 5.33707e-19
cc_8 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.00168612f
cc_9 N_VSS_XI0.X0_PGD N_VDD_XI3.X0_PGD 0.00189944f
cc_10 N_VSS_XI5.X0_PGD N_VDD_XI4.X0_PGD 0.00180681f
cc_11 N_VSS_c_11_p N_VDD_c_152_n 0.00168612f
cc_12 N_VSS_c_12_p N_VDD_c_153_n 0.00189944f
cc_13 N_VSS_c_13_p N_VDD_c_154_n 0.00180681f
cc_14 N_VSS_XI1.X0_S N_VDD_c_155_n 9.5668e-19
cc_15 N_VSS_c_15_p N_VDD_c_155_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_155_n 0.00321182f
cc_17 N_VSS_c_17_p N_VDD_c_155_n 0.00182807f
cc_18 N_VSS_c_15_p N_VDD_c_159_n 5.16845e-19
cc_19 N_VSS_c_3_p N_VDD_c_159_n 2.61925e-19
cc_20 N_VSS_c_20_p N_VDD_c_159_n 4.48125e-19
cc_21 N_VSS_c_7_p N_VDD_c_159_n 0.00922264f
cc_22 N_VSS_c_22_p N_VDD_c_163_n 0.00105444f
cc_23 N_VSS_c_23_p N_VDD_c_164_n 0.00239254f
cc_24 N_VSS_c_4_p N_VDD_c_164_n 9.55109e-19
cc_25 N_VSS_c_13_p N_VDD_c_166_n 2.43144e-19
cc_26 N_VSS_c_23_p N_VDD_c_166_n 0.00161703f
cc_27 N_VSS_c_4_p N_VDD_c_166_n 2.03837e-19
cc_28 N_VSS_c_7_p N_VDD_c_166_n 0.00131925f
cc_29 N_VSS_c_29_p N_VDD_c_166_n 0.00399563f
cc_30 N_VSS_c_30_p N_VDD_c_166_n 7.74609e-19
cc_31 N_VSS_c_3_p N_VDD_c_172_n 0.00179177f
cc_32 N_VSS_c_32_p N_VDD_c_172_n 3.92901e-19
cc_33 N_VSS_c_33_p N_VDD_c_172_n 8.51944e-19
cc_34 N_VSS_c_34_p N_VDD_c_172_n 3.99794e-19
cc_35 N_VSS_c_12_p N_VDD_c_176_n 3.37151e-19
cc_36 N_VSS_c_33_p N_VDD_c_176_n 0.00141228f
cc_37 N_VSS_c_34_p N_VDD_c_176_n 0.00112249f
cc_38 N_VSS_c_38_p N_VDD_c_176_n 0.00402042f
cc_39 N_VSS_c_39_p N_VDD_c_176_n 0.00326829f
cc_40 N_VSS_c_40_p N_VDD_c_176_n 7.74609e-19
cc_41 N_VSS_c_38_p N_VDD_c_182_n 0.00142104f
cc_42 N_VSS_c_23_p N_VDD_c_183_n 9.29543e-19
cc_43 N_VSS_c_4_p N_VDD_c_183_n 3.82294e-19
cc_44 N_VSS_XI4.X0_S N_VDD_c_185_n 3.7884e-19
cc_45 N_VSS_c_45_p N_VDD_c_185_n 4.73473e-19
cc_46 N_VSS_c_29_p N_VDD_c_185_n 0.00432522f
cc_47 N_VSS_c_45_p N_VDD_c_188_n 2.14355e-19
cc_48 N_VSS_c_48_p N_VDD_c_188_n 5.52785e-19
cc_49 N_VSS_XI4.X0_S N_VDD_c_190_n 9.5668e-19
cc_50 N_VSS_c_45_p N_VDD_c_190_n 0.00165395f
cc_51 N_VSS_c_51_p N_VDD_c_190_n 0.00302432f
cc_52 N_VSS_c_52_p N_VDD_c_190_n 0.00617602f
cc_53 N_VSS_c_53_p N_VDD_c_190_n 8.91588e-19
cc_54 N_VSS_c_33_p N_VDD_c_195_n 4.43871e-19
cc_55 N_VSS_c_34_p N_VDD_c_195_n 3.66936e-19
cc_56 N_VSS_c_39_p N_VDD_c_195_n 0.00106633f
cc_57 N_VSS_c_52_p N_VDD_c_195_n 0.00303537f
cc_58 N_VSS_c_3_p N_VDD_c_199_n 6.19689e-19
cc_59 N_VSS_c_20_p N_VDD_c_199_n 3.8721e-19
cc_60 N_VSS_c_15_p N_VDD_c_201_n 0.00303908f
cc_61 N_VSS_c_7_p N_VDD_c_201_n 2.94014e-19
cc_62 N_VSS_c_7_p N_VDD_c_203_n 0.00116322f
cc_63 N_VSS_c_29_p N_VDD_c_204_n 0.00102846f
cc_64 N_VSS_c_52_p N_VDD_c_205_n 0.00116512f
cc_65 N_VSS_c_3_p N_VDD_c_206_n 3.86162e-19
cc_66 N_VSS_c_20_p N_VDD_c_206_n 6.0892e-19
cc_67 N_VSS_c_3_p N_VDD_c_208_n 5.29489e-19
cc_68 N_VSS_c_33_p N_VDD_c_208_n 3.48267e-19
cc_69 N_VSS_c_34_p N_VDD_c_208_n 8.07896e-19
cc_70 N_VSS_c_23_p N_VDD_c_211_n 3.48267e-19
cc_71 N_VSS_c_4_p N_VDD_c_211_n 8.0279e-19
cc_72 N_VSS_XI1.X0_S N_CKN_XI1.X0_D 3.43419e-19
cc_73 N_VSS_c_15_p N_CKN_XI1.X0_D 3.48267e-19
cc_74 N_VSS_XI1.X0_S N_CKN_c_268_n 3.48267e-19
cc_75 N_VSS_c_15_p N_CKN_c_268_n 0.00105962f
cc_76 N_VSS_c_3_p N_CKN_c_268_n 7.53164e-19
cc_77 N_VSS_c_7_p N_CKN_c_268_n 5.38016e-19
cc_78 N_VSS_c_29_p N_CKN_c_272_n 2.21217e-19
cc_79 N_VSS_c_52_p N_CKN_c_272_n 0.00111539f
cc_80 N_VSS_c_3_p N_CKN_c_274_n 0.00220607f
cc_81 N_VSS_c_32_p N_CKN_c_274_n 8.60018e-19
cc_82 N_VSS_c_23_p N_CKN_c_274_n 2.36534e-19
cc_83 N_VSS_c_33_p N_CKN_c_274_n 7.62758e-19
cc_84 N_VSS_c_7_p N_CKN_c_274_n 0.00158805f
cc_85 N_VSS_c_85_p N_CKN_c_274_n 8.14378e-19
cc_86 N_VSS_c_38_p N_CKN_c_274_n 9.16986e-19
cc_87 N_VSS_c_29_p N_CKN_c_274_n 0.00110784f
cc_88 N_VSS_c_4_p N_D_XI5.X0_CG 0.00265616f
cc_89 N_VSS_c_89_p N_D_c_305_n 9.49637e-19
cc_90 N_VSS_XI5.X0_PGD N_D_c_306_n 3.8966e-19
cc_91 N_VSS_XI0.X0_PGD N_D_c_306_n 2.22031e-19
cc_92 N_VSS_c_3_p N_D_c_308_n 6.13924e-19
cc_93 N_VSS_c_23_p N_D_c_308_n 5.5494e-19
cc_94 N_VSS_c_20_p N_D_c_308_n 3.48267e-19
cc_95 N_VSS_c_4_p N_D_c_308_n 4.56568e-19
cc_96 N_VSS_c_3_p N_D_c_312_n 3.48267e-19
cc_97 N_VSS_c_23_p N_D_c_312_n 4.56568e-19
cc_98 N_VSS_c_20_p N_D_c_312_n 6.88619e-19
cc_99 N_VSS_c_4_p N_D_c_312_n 6.1245e-19
cc_100 N_VSS_XI4.X0_S N_X_XI5.X0_D 3.43419e-19
cc_101 N_VSS_c_45_p N_X_XI5.X0_D 3.48267e-19
cc_102 N_VSS_c_34_p N_X_XI0.X0_CG 0.00105235f
cc_103 N_VSS_XI5.X0_PGD N_X_c_334_n 2.09879e-19
cc_104 N_VSS_XI0.X0_PGD N_X_c_334_n 3.99472e-19
cc_105 N_VSS_c_38_p N_X_c_336_n 2.5064e-19
cc_106 N_VSS_XI4.X0_S N_X_c_337_n 3.48267e-19
cc_107 N_VSS_c_3_p N_X_c_337_n 4.71026e-19
cc_108 N_VSS_c_45_p N_X_c_337_n 5.69026e-19
cc_109 N_VSS_c_52_p N_X_c_337_n 2.04792e-19
cc_110 N_VSS_c_3_p N_X_c_341_n 0.00157847f
cc_111 N_VSS_c_52_p N_X_c_341_n 3.24972e-19
cc_112 N_VSS_c_3_p N_X_c_343_n 3.48267e-19
cc_113 N_VSS_c_4_p N_X_c_343_n 2.00604e-19
cc_114 N_VSS_XI3.X0_S N_Q_XI3.X0_D 3.43419e-19
cc_115 N_VSS_c_32_p N_Q_XI3.X0_D 3.48267e-19
cc_116 N_VSS_XI3.X0_S Q 3.48267e-19
cc_117 N_VSS_c_32_p Q 4.99861e-19
cc_118 N_CK_c_122_n N_VDD_XI1.X0_PGD 4.16623e-19
cc_119 N_CK_XI5.X0_PGS N_VDD_XI4.X0_PGD 2.40707e-19
cc_120 N_CK_c_123_n N_VDD_c_154_n 2.40707e-19
cc_121 CK N_VDD_c_155_n 5.04211e-19
cc_122 N_CK_c_129_p N_VDD_c_155_n 5.23418e-19
cc_123 N_CK_c_122_n N_VDD_c_159_n 0.00141086f
cc_124 CK N_VDD_c_159_n 0.00141439f
cc_125 N_CK_c_129_p N_VDD_c_159_n 0.00120361f
cc_126 N_CK_XI5.X0_PGS N_VDD_c_164_n 2.38687e-19
cc_127 N_CK_c_123_n N_VDD_c_164_n 5.38952e-19
cc_128 CK N_VDD_c_164_n 3.91916e-19
cc_129 N_CK_c_129_p N_VDD_c_164_n 2.80271e-19
cc_130 CK N_VDD_c_199_n 6.07878e-19
cc_131 N_CK_c_129_p N_VDD_c_199_n 4.67029e-19
cc_132 CK N_VDD_c_206_n 4.56568e-19
cc_133 N_CK_c_129_p N_VDD_c_206_n 0.00211811f
cc_134 N_CK_XI5.X0_PGS N_CKN_XI4.X0_PGS 4.11563e-19
cc_135 N_CK_XI5.X0_PGS N_CKN_c_283_n 2.73384e-19
cc_136 N_CK_XI5.X0_PGS N_D_XI5.X0_CG 4.28946e-19
cc_137 N_CK_XI5.X0_PGS N_D_XI4.X0_CG 2.59344e-19
cc_138 N_CK_XI5.X0_PGS N_D_c_312_n 0.00300565f
cc_139 N_CK_XI5.X0_PGS N_X_XI0.X0_CG 2.6404e-19
cc_140 N_CK_XI5.X0_PGS N_X_c_346_n 4.97357e-19
cc_141 N_CK_XI5.X0_PGS N_X_c_343_n 0.00630896f
cc_142 N_VDD_XI2.X0_S N_CKN_XI1.X0_D 3.43419e-19
cc_143 N_VDD_c_190_n N_CKN_XI4.X0_PGS 5.54393e-19
cc_144 N_VDD_c_190_n N_CKN_c_283_n 8.21431e-19
cc_145 N_VDD_XI2.X0_S N_CKN_c_268_n 3.48267e-19
cc_146 N_VDD_c_159_n N_CKN_c_268_n 5.01863e-19
cc_147 N_VDD_c_164_n N_CKN_c_268_n 5.35331e-19
cc_148 N_VDD_c_199_n N_CKN_c_268_n 6.42405e-19
cc_149 N_VDD_c_190_n N_CKN_c_272_n 7.71262e-19
cc_150 N_VDD_c_159_n N_CKN_c_274_n 4.68667e-19
cc_151 N_VDD_c_166_n N_CKN_c_274_n 3.15582e-19
cc_152 N_VDD_c_176_n N_CKN_c_274_n 4.71809e-19
cc_153 N_VDD_c_183_n N_CKN_c_274_n 2.56401e-19
cc_154 N_VDD_c_211_n N_D_XI4.X0_CG 0.00105644f
cc_155 N_VDD_XI3.X0_PGD N_D_c_306_n 2.08865e-19
cc_156 N_VDD_XI4.X0_PGD N_D_c_306_n 4.04053e-19
cc_157 N_VDD_XI2.X0_S N_X_XI5.X0_D 3.43419e-19
cc_158 N_VDD_c_164_n N_X_XI5.X0_D 3.48267e-19
cc_159 N_VDD_c_166_n N_X_XI5.X0_D 3.7884e-19
cc_160 N_VDD_c_208_n N_X_c_346_n 0.00269538f
cc_161 N_VDD_XI3.X0_PGD N_X_c_334_n 3.93054e-19
cc_162 N_VDD_XI4.X0_PGD N_X_c_334_n 2.22031e-19
cc_163 N_VDD_c_250_p N_X_c_354_n 8.95961e-19
cc_164 N_VDD_c_208_n N_X_c_354_n 2.97161e-19
cc_165 N_VDD_XI2.X0_S N_X_c_337_n 3.48267e-19
cc_166 N_VDD_c_164_n N_X_c_337_n 6.883e-19
cc_167 N_VDD_c_166_n N_X_c_337_n 5.3319e-19
cc_168 N_VDD_c_190_n N_X_c_337_n 8.74231e-19
cc_169 N_VDD_c_172_n N_X_c_341_n 6.5515e-19
cc_170 N_VDD_c_208_n N_X_c_341_n 4.80549e-19
cc_171 N_VDD_c_172_n N_X_c_343_n 4.85469e-19
cc_172 N_VDD_c_208_n N_X_c_343_n 6.1245e-19
cc_173 N_VDD_XI0.X0_S N_Q_XI3.X0_D 3.43419e-19
cc_174 N_VDD_c_176_n N_Q_XI3.X0_D 3.7884e-19
cc_175 N_VDD_c_188_n N_Q_XI3.X0_D 3.72199e-19
cc_176 N_VDD_XI0.X0_S Q 3.48267e-19
cc_177 N_VDD_c_176_n Q 5.12447e-19
cc_178 N_VDD_c_188_n Q 7.06537e-19
cc_179 N_CKN_XI4.X0_PGS N_D_XI4.X0_CG 0.00392964f
cc_180 N_CKN_XI4.X0_PGS N_X_c_334_n 0.00402435f
cc_181 N_CKN_c_283_n N_X_c_336_n 5.71169e-19
cc_182 N_CKN_c_274_n N_X_c_336_n 0.00120349f
cc_183 N_CKN_c_268_n N_X_c_337_n 2.66307e-19
cc_184 N_CKN_c_272_n N_X_c_337_n 8.08281e-19
cc_185 N_CKN_c_274_n N_X_c_337_n 6.2695e-19
cc_186 N_CKN_c_274_n N_X_c_341_n 7.98434e-19
cc_187 N_D_c_306_n N_X_c_334_n 0.00454934f
cc_188 N_D_c_306_n N_X_c_337_n 2.96904e-19
cc_189 N_D_c_308_n N_X_c_337_n 0.00151915f
cc_190 N_D_c_312_n N_X_c_337_n 9.22925e-19
cc_191 N_D_c_308_n N_X_c_341_n 0.00146206f
cc_192 N_D_c_312_n N_X_c_341_n 0.00103457f
cc_193 N_D_c_308_n N_X_c_343_n 4.56568e-19
cc_194 N_D_c_312_n N_X_c_343_n 0.00373298f
cc_195 N_X_c_336_n N_Q_XI3.X0_D 5.75967e-19
cc_196 N_X_c_336_n Q 8.57825e-19
*
.ends
*
*
.subckt DFFQ1_HPNW4 CK D Q VDD VSS
xgate (VSS CK VDD D Q) G3_DFFQ1_N1_2
.ends
*
* File: G1_INV1_N1.pex.netlist
* Created: Fri Feb 18 12:29:10 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*




.subckt G1_INV1_N1_2 VDD A VSS Z
*
* Z	Z
* VSS	VSS
* A	A
* VDD	VDD
XI2.X0 N_Z_XI2.X0_D N_VSS_XI2.X0_PGD N_A_XI2.X0_CG N_VSS_XI2.X0_PGD
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI1.X0 N_Z_XI2.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW4
*
x_PM_G1_INV1_N1_VDD N_VDD_XI2.X0_S N_VDD_XI1.X0_PGD N_VDD_c_5_p N_VDD_c_4_p
+ N_VDD_c_6_p N_VDD_c_9_p VDD N_VDD_c_1_p Vss PM_G1_INV1_N1_VDD
x_PM_G1_INV1_N1_A N_A_XI2.X0_CG N_A_XI1.X0_CG N_A_c_29_p N_A_c_25_n A N_A_c_27_p
+ N_A_c_28_p Vss PM_G1_INV1_N1_A
x_PM_G1_INV1_N1_VSS N_VSS_XI2.X0_PGD N_VSS_XI1.X0_S N_VSS_c_34_n N_VSS_c_36_n
+ N_VSS_c_40_n N_VSS_c_42_n N_VSS_c_45_n N_VSS_c_46_n VSS Vss PM_G1_INV1_N1_VSS
x_PM_G1_INV1_N1_Z N_Z_XI2.X0_D Z Vss PM_G1_INV1_N1_Z
cc_1 N_VDD_c_1_p N_A_XI1.X0_CG 8.21222e-19
cc_2 N_VDD_XI1.X0_PGD N_A_c_25_n 4.26524e-19
cc_3 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00171093f
cc_4 N_VDD_c_4_p N_VSS_XI2.X0_PGD 4.197e-19
cc_5 N_VDD_c_5_p N_VSS_c_34_n 0.00171093f
cc_6 N_VDD_c_6_p N_VSS_c_34_n 4.82774e-19
cc_7 N_VDD_c_4_p N_VSS_c_36_n 0.00304634f
cc_8 N_VDD_c_6_p N_VSS_c_36_n 0.0015849f
cc_9 N_VDD_c_9_p N_VSS_c_36_n 9.51078e-19
cc_10 N_VDD_c_1_p N_VSS_c_36_n 3.5189e-19
cc_11 N_VDD_c_4_p N_VSS_c_40_n 3.08259e-19
cc_12 N_VDD_c_9_p N_VSS_c_40_n 0.00107037f
cc_13 N_VDD_c_4_p N_VSS_c_42_n 9.54992e-19
cc_14 N_VDD_c_9_p N_VSS_c_42_n 3.83199e-19
cc_15 N_VDD_c_1_p N_VSS_c_42_n 7.7548e-19
cc_16 N_VDD_c_6_p N_VSS_c_45_n 0.005791f
cc_17 N_VDD_c_6_p N_VSS_c_46_n 0.00172748f
cc_18 N_VDD_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_19 N_VDD_c_4_p N_Z_XI2.X0_D 3.48267e-19
cc_20 N_VDD_c_6_p N_Z_XI2.X0_D 3.55567e-19
cc_21 N_VDD_XI2.X0_S Z 3.48267e-19
cc_22 N_VDD_c_4_p Z 7.06424e-19
cc_23 N_VDD_c_6_p Z 4.789e-19
cc_24 N_A_c_25_n N_VSS_XI2.X0_PGD 4.21166e-19
cc_25 N_A_c_27_p N_VSS_c_36_n 0.00103813f
cc_26 N_A_c_28_p N_VSS_c_36_n 4.99367e-19
cc_27 N_A_c_29_p N_VSS_c_42_n 0.00250475f
cc_28 N_A_c_27_p N_VSS_c_42_n 4.99367e-19
cc_29 N_A_c_28_p N_VSS_c_42_n 0.0014909f
cc_30 N_VSS_XI1.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_31 N_VSS_c_40_n N_Z_XI2.X0_D 3.48267e-19
cc_32 N_VSS_XI1.X0_S Z 3.48267e-19
cc_33 N_VSS_c_40_n Z 7.85754e-19
cc_34 N_VSS_c_45_n Z 2.54816e-19
*
.ends
*
*
.subckt INV1_HPNW4 A Y VDD VSS
xgate (VDD A VSS Y) G1_INV1_N1_2
.ends
*
* File: G3_LATQ1_N1.pex.netlist
* Created: Tue Apr  5 11:43:13 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*







.subckt G3_LATQ1_N1_2 VDD VSS G Q D
*
* D	D
* Q	Q
* G	G
* VSS	VSS
* VDD	VDD
XI2.X0 N_GN_XI2.X0_D N_VSS_XI2.X0_PGD N_G_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI0.X0 N_Q_XI0.X0_D N_VDD_XI0.X0_PGD N_QN_XI0.X0_CG N_VDD_XI0.X0_PGS
+ N_VSS_XI0.X0_S TIGFET_HPNW4
XI1.X0 N_GN_XI2.X0_D N_VDD_XI1.X0_PGD N_G_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI3.X0 N_Q_XI0.X0_D N_VSS_XI3.X0_PGD N_QN_XI3.X0_CG N_VSS_XI3.X0_PGS
+ N_VDD_XI3.X0_S TIGFET_HPNW4
XI5.X0 N_QN_XI5.X0_D N_VDD_XI5.X0_PGD N_D_XI5.X0_CG N_G_XI5.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI4.X0 N_QN_XI4.X0_D N_VSS_XI4.X0_PGD N_D_XI4.X0_CG N_GN_XI4.X0_PGS
+ N_VDD_XI3.X0_S TIGFET_HPNW4
*
x_PM_G3_LATQ1_N1_VDD N_VDD_XI2.X0_S N_VDD_XI0.X0_PGD N_VDD_XI0.X0_PGS
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI3.X0_S N_VDD_XI5.X0_PGD N_VDD_c_10_p
+ N_VDD_c_58_p N_VDD_c_7_p N_VDD_c_47_p N_VDD_c_16_p N_VDD_c_3_p N_VDD_c_8_p
+ N_VDD_c_38_p N_VDD_c_14_p N_VDD_c_15_p N_VDD_c_42_p N_VDD_c_20_p N_VDD_c_11_p
+ N_VDD_c_18_p N_VDD_c_5_p N_VDD_c_35_p N_VDD_c_41_p VDD N_VDD_c_23_p
+ N_VDD_c_19_p Vss PM_G3_LATQ1_N1_VDD
x_PM_G3_LATQ1_N1_VSS N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS N_VSS_XI0.X0_S
+ N_VSS_XI1.X0_S N_VSS_XI3.X0_PGD N_VSS_XI3.X0_PGS N_VSS_XI4.X0_PGD N_VSS_c_98_n
+ N_VSS_c_100_n N_VSS_c_101_n N_VSS_c_103_n N_VSS_c_104_n N_VSS_c_107_n
+ N_VSS_c_111_n N_VSS_c_115_n N_VSS_c_116_n N_VSS_c_120_n N_VSS_c_124_n
+ N_VSS_c_127_n N_VSS_c_128_n N_VSS_c_129_n N_VSS_c_130_n N_VSS_c_133_n
+ N_VSS_c_134_n N_VSS_c_135_n N_VSS_c_136_n VSS Vss PM_G3_LATQ1_N1_VSS
x_PM_G3_LATQ1_N1_G N_G_XI2.X0_CG N_G_XI1.X0_CG N_G_XI5.X0_PGS N_G_c_183_n
+ N_G_c_177_n N_G_c_179_n G N_G_c_181_n Vss PM_G3_LATQ1_N1_G
x_PM_G3_LATQ1_N1_QN N_QN_XI0.X0_CG N_QN_XI3.X0_CG N_QN_XI5.X0_D N_QN_XI4.X0_D
+ N_QN_c_205_n N_QN_c_206_n N_QN_c_208_n N_QN_c_210_n N_QN_c_213_n N_QN_c_215_n
+ N_QN_c_218_n N_QN_c_221_n Vss PM_G3_LATQ1_N1_QN
x_PM_G3_LATQ1_N1_GN N_GN_XI2.X0_D N_GN_XI4.X0_PGS N_GN_c_254_n N_GN_c_256_n
+ N_GN_c_279_n N_GN_c_285_n N_GN_c_260_n N_GN_c_262_n Vss PM_G3_LATQ1_N1_GN
x_PM_G3_LATQ1_N1_Q N_Q_XI0.X0_D Q Vss PM_G3_LATQ1_N1_Q
x_PM_G3_LATQ1_N1_D N_D_XI5.X0_CG N_D_XI4.X0_CG N_D_c_314_n D Vss
+ PM_G3_LATQ1_N1_D
cc_1 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00175469f
cc_2 N_VDD_XI0.X0_PGS N_VSS_XI2.X0_PGS 2.27468e-19
cc_3 N_VDD_c_3_p N_VSS_XI0.X0_S 9.5668e-19
cc_4 N_VDD_XI0.X0_PGD N_VSS_XI3.X0_PGD 0.00173629f
cc_5 N_VDD_c_5_p N_VSS_XI3.X0_PGS 2.46127e-19
cc_6 N_VDD_XI5.X0_PGD N_VSS_XI4.X0_PGD 2.27468e-19
cc_7 N_VDD_c_7_p N_VSS_c_98_n 0.00175469f
cc_8 N_VDD_c_8_p N_VSS_c_98_n 3.60588e-19
cc_9 N_VDD_c_8_p N_VSS_c_100_n 3.60588e-19
cc_10 N_VDD_c_10_p N_VSS_c_101_n 0.00173629f
cc_11 N_VDD_c_11_p N_VSS_c_101_n 2.60334e-19
cc_12 N_VDD_c_5_p N_VSS_c_103_n 7.75484e-19
cc_13 N_VDD_c_3_p N_VSS_c_104_n 0.00165395f
cc_14 N_VDD_c_14_p N_VSS_c_104_n 7.6714e-19
cc_15 N_VDD_c_15_p N_VSS_c_104_n 5.16845e-19
cc_16 N_VDD_c_16_p N_VSS_c_107_n 4.43871e-19
cc_17 N_VDD_c_8_p N_VSS_c_107_n 0.00161703f
cc_18 N_VDD_c_18_p N_VSS_c_107_n 9.31718e-19
cc_19 N_VDD_c_19_p N_VSS_c_107_n 3.48267e-19
cc_20 N_VDD_c_20_p N_VSS_c_111_n 9.36729e-19
cc_21 N_VDD_c_11_p N_VSS_c_111_n 0.00141228f
cc_22 N_VDD_c_5_p N_VSS_c_111_n 0.00291977f
cc_23 N_VDD_c_23_p N_VSS_c_111_n 3.5189e-19
cc_24 N_VDD_c_18_p N_VSS_c_115_n 0.00102583f
cc_25 N_VDD_c_16_p N_VSS_c_116_n 3.66936e-19
cc_26 N_VDD_c_8_p N_VSS_c_116_n 2.03837e-19
cc_27 N_VDD_c_18_p N_VSS_c_116_n 3.99794e-19
cc_28 N_VDD_c_19_p N_VSS_c_116_n 8.07896e-19
cc_29 N_VDD_c_20_p N_VSS_c_120_n 3.86045e-19
cc_30 N_VDD_c_11_p N_VSS_c_120_n 0.00112249f
cc_31 N_VDD_c_5_p N_VSS_c_120_n 9.54992e-19
cc_32 N_VDD_c_23_p N_VSS_c_120_n 8.1718e-19
cc_33 N_VDD_c_16_p N_VSS_c_124_n 0.00303537f
cc_34 N_VDD_c_3_p N_VSS_c_124_n 0.00544275f
cc_35 N_VDD_c_35_p N_VSS_c_124_n 0.00116512f
cc_36 N_VDD_c_3_p N_VSS_c_127_n 0.00305967f
cc_37 N_VDD_c_8_p N_VSS_c_128_n 0.00343927f
cc_38 N_VDD_c_38_p N_VSS_c_129_n 0.00106317f
cc_39 N_VDD_c_15_p N_VSS_c_130_n 0.00355199f
cc_40 N_VDD_c_11_p N_VSS_c_130_n 0.00567045f
cc_41 N_VDD_c_41_p N_VSS_c_130_n 9.48532e-19
cc_42 N_VDD_c_42_p N_VSS_c_133_n 0.00105938f
cc_43 N_VDD_c_8_p N_VSS_c_134_n 0.00557463f
cc_44 N_VDD_c_3_p N_VSS_c_135_n 8.91588e-19
cc_45 N_VDD_c_8_p N_VSS_c_136_n 7.74609e-19
cc_46 N_VDD_c_19_p N_G_XI1.X0_CG 8.09841e-19
cc_47 N_VDD_c_47_p N_G_XI5.X0_PGS 0.00162079f
cc_48 N_VDD_XI0.X0_PGD N_G_c_177_n 2.22031e-19
cc_49 N_VDD_XI1.X0_PGD N_G_c_177_n 3.93641e-19
cc_50 N_VDD_XI1.X0_PGS N_G_c_179_n 4.05198e-19
cc_51 N_VDD_c_3_p G 3.46645e-19
cc_52 N_VDD_c_3_p N_G_c_181_n 4.43544e-19
cc_53 N_VDD_XI3.X0_S N_QN_XI4.X0_D 3.43419e-19
cc_54 N_VDD_c_5_p N_QN_XI4.X0_D 3.48267e-19
cc_55 N_VDD_c_23_p N_QN_c_205_n 0.00269246f
cc_56 N_VDD_XI0.X0_PGD N_QN_c_206_n 4.05198e-19
cc_57 N_VDD_XI1.X0_PGD N_QN_c_206_n 2.0936e-19
cc_58 N_VDD_c_58_p N_QN_c_208_n 9.69462e-19
cc_59 N_VDD_c_23_p N_QN_c_208_n 2.60536e-19
cc_60 N_VDD_c_3_p N_QN_c_210_n 4.49462e-19
cc_61 N_VDD_c_20_p N_QN_c_210_n 4.57093e-19
cc_62 N_VDD_c_23_p N_QN_c_210_n 4.4444e-19
cc_63 N_VDD_XI3.X0_S N_QN_c_213_n 3.48267e-19
cc_64 N_VDD_c_5_p N_QN_c_213_n 9.00822e-19
cc_65 N_VDD_c_8_p N_QN_c_215_n 4.48879e-19
cc_66 N_VDD_c_11_p N_QN_c_215_n 3.93728e-19
cc_67 N_VDD_c_5_p N_QN_c_215_n 3.58217e-19
cc_68 N_VDD_c_3_p N_QN_c_218_n 6.61926e-19
cc_69 N_VDD_c_20_p N_QN_c_218_n 4.85469e-19
cc_70 N_VDD_c_23_p N_QN_c_218_n 6.1245e-19
cc_71 N_VDD_c_3_p N_QN_c_221_n 4.64547e-19
cc_72 N_VDD_XI2.X0_S N_GN_XI2.X0_D 3.43419e-19
cc_73 N_VDD_c_8_p N_GN_XI2.X0_D 3.7884e-19
cc_74 N_VDD_c_14_p N_GN_XI2.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_PGS N_GN_c_254_n 3.40151e-19
cc_76 N_VDD_c_47_p N_GN_c_254_n 3.20239e-19
cc_77 N_VDD_XI2.X0_S N_GN_c_256_n 3.48267e-19
cc_78 N_VDD_c_3_p N_GN_c_256_n 6.12365e-19
cc_79 N_VDD_c_8_p N_GN_c_256_n 5.32769e-19
cc_80 N_VDD_c_14_p N_GN_c_256_n 7.89245e-19
cc_81 N_VDD_c_18_p N_GN_c_260_n 2.2082e-19
cc_82 N_VDD_c_19_p N_GN_c_260_n 2.46105e-19
cc_83 N_VDD_c_18_p N_GN_c_262_n 2.68489e-19
cc_84 N_VDD_c_19_p N_GN_c_262_n 5.71759e-19
cc_85 N_VDD_XI3.X0_S N_Q_XI0.X0_D 3.43419e-19
cc_86 N_VDD_c_11_p N_Q_XI0.X0_D 3.7884e-19
cc_87 N_VDD_c_5_p N_Q_XI0.X0_D 3.48267e-19
cc_88 N_VDD_XI3.X0_S Q 3.48267e-19
cc_89 N_VDD_c_11_p Q 5.12447e-19
cc_90 N_VDD_c_5_p Q 7.06424e-19
cc_91 N_VDD_c_47_p N_D_XI5.X0_CG 4.07085e-19
cc_92 N_VSS_c_116_n N_G_XI2.X0_CG 0.00265616f
cc_93 N_VSS_c_116_n N_G_c_183_n 9.49637e-19
cc_94 N_VSS_XI2.X0_PGD N_G_c_177_n 3.99472e-19
cc_95 N_VSS_XI3.X0_PGD N_G_c_177_n 2.0936e-19
cc_96 N_VSS_c_107_n G 5.5494e-19
cc_97 N_VSS_c_116_n G 4.56568e-19
cc_98 N_VSS_c_124_n G 3.38887e-19
cc_99 N_VSS_c_107_n N_G_c_181_n 4.56568e-19
cc_100 N_VSS_c_116_n N_G_c_181_n 6.1245e-19
cc_101 N_VSS_c_120_n N_QN_XI3.X0_CG 8.05748e-19
cc_102 N_VSS_XI1.X0_S N_QN_XI5.X0_D 3.43419e-19
cc_103 N_VSS_c_115_n N_QN_XI5.X0_D 3.48267e-19
cc_104 N_VSS_XI2.X0_PGD N_QN_c_206_n 2.22031e-19
cc_105 N_VSS_XI3.X0_PGD N_QN_c_206_n 3.89061e-19
cc_106 N_VSS_c_130_n N_QN_c_210_n 2.91026e-19
cc_107 N_VSS_c_115_n N_QN_c_213_n 8.97415e-19
cc_108 N_VSS_c_111_n N_QN_c_215_n 3.5258e-19
cc_109 N_VSS_c_115_n N_QN_c_215_n 7.99552e-19
cc_110 N_VSS_c_130_n N_QN_c_215_n 6.85871e-19
cc_111 N_VSS_c_134_n N_QN_c_215_n 9.55516e-19
cc_112 N_VSS_c_107_n N_QN_c_221_n 5.43247e-19
cc_113 N_VSS_c_124_n N_QN_c_221_n 0.00168288f
cc_114 N_VSS_XI1.X0_S N_GN_XI2.X0_D 3.43419e-19
cc_115 N_VSS_c_115_n N_GN_XI2.X0_D 3.48267e-19
cc_116 N_VSS_c_103_n N_GN_XI4.X0_PGS 0.00163489f
cc_117 N_VSS_XI3.X0_PGS N_GN_c_254_n 6.77138e-19
cc_118 N_VSS_c_103_n N_GN_c_254_n 2.57527e-19
cc_119 N_VSS_XI1.X0_S N_GN_c_256_n 3.48267e-19
cc_120 N_VSS_c_115_n N_GN_c_256_n 4.97497e-19
cc_121 N_VSS_c_124_n N_GN_c_256_n 4.46497e-19
cc_122 N_VSS_c_120_n N_GN_c_260_n 2.46105e-19
cc_123 N_VSS_c_111_n N_GN_c_262_n 2.52506e-19
cc_124 N_VSS_c_120_n N_GN_c_262_n 5.99566e-19
cc_125 N_VSS_XI0.X0_S N_Q_XI0.X0_D 3.43419e-19
cc_126 N_VSS_c_104_n N_Q_XI0.X0_D 3.48267e-19
cc_127 N_VSS_XI0.X0_S Q 3.48267e-19
cc_128 N_VSS_c_104_n Q 7.78122e-19
cc_129 N_VSS_c_103_n N_D_XI5.X0_CG 4.07085e-19
cc_130 N_G_c_177_n N_QN_c_206_n 0.003965f
cc_131 G N_QN_c_210_n 5.07332e-19
cc_132 N_G_c_181_n N_QN_c_210_n 4.54925e-19
cc_133 N_G_c_181_n N_QN_c_218_n 0.00269321f
cc_134 N_G_c_179_n N_GN_c_254_n 0.00851239f
cc_135 N_G_c_177_n N_GN_c_256_n 3.2445e-19
cc_136 G N_GN_c_256_n 0.00153131f
cc_137 N_G_c_181_n N_GN_c_256_n 9.18093e-19
cc_138 N_G_c_177_n N_GN_c_279_n 3.7133e-19
cc_139 N_G_c_177_n N_GN_c_262_n 9.94034e-19
cc_140 N_G_c_181_n N_GN_c_262_n 2.41671e-19
cc_141 N_G_XI5.X0_PGS N_D_XI5.X0_CG 0.00409312f
cc_142 N_QN_c_206_n N_GN_XI4.X0_PGS 0.00182388f
cc_143 N_QN_c_213_n N_GN_c_256_n 7.80248e-19
cc_144 N_QN_c_215_n N_GN_c_279_n 8.96813e-19
cc_145 N_QN_c_215_n N_GN_c_285_n 0.00118168f
cc_146 N_QN_c_215_n N_GN_c_260_n 9.24681e-19
cc_147 N_QN_c_206_n N_GN_c_262_n 8.57779e-19
cc_148 N_QN_c_218_n N_GN_c_262_n 2.75519e-19
cc_149 N_QN_c_206_n N_D_XI5.X0_CG 3.26559e-19
cc_150 N_QN_c_213_n N_D_XI5.X0_CG 0.00101289f
cc_151 N_QN_c_213_n N_D_c_314_n 0.00127983f
cc_152 N_QN_c_213_n D 0.00141415f
cc_153 N_QN_c_215_n D 0.00146947f
cc_154 N_GN_c_285_n N_Q_XI0.X0_D 5.19956e-19
cc_155 N_GN_c_285_n Q 6.79271e-19
cc_156 N_GN_XI4.X0_PGS N_D_XI5.X0_CG 0.00503657f
cc_157 N_GN_c_254_n N_D_c_314_n 0.00333193f
cc_158 N_GN_c_260_n N_D_c_314_n 3.73302e-19
cc_159 N_GN_c_262_n N_D_c_314_n 8.5422e-19
cc_160 N_GN_c_260_n D 2.88184e-19
cc_161 N_GN_c_262_n D 3.48267e-19
*
.ends
*
*
.subckt LATQ1_HPNW4 D G Q VDD VSS
xgate (VDD VSS G Q D) G3_LATQ1_N1_2
.ends
*
* File: G4_MAJ3_N1.pex.netlist
* Created: Wed Mar  2 17:07:12 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*








.subckt G4_MAJ3_N1_2 VDD VSS A B C Z
*
* Z	Z
* C	C
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI6.X0 N_BI_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW4
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI5.X0 N_VSS_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_BI_XI6.X0_D TIGFET_HPNW4
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW4
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_BI_XI2.X0_CG N_AI_XI2.X0_PGD N_A_XI2.X0_S
+ TIGFET_HPNW4
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_B_XI4.X0_CG N_AI_XI4.X0_PGD N_C_XI4.X0_S
+ TIGFET_HPNW4
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_B_XI3.X0_CG N_A_XI3.X0_PGD N_A_XI3.X0_S
+ TIGFET_HPNW4
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_BI_XI1.X0_CG N_A_XI1.X0_PGD N_C_XI1.X0_S
+ TIGFET_HPNW4
*
x_PM_G4_MAJ3_N1_VDD N_VDD_XI6.X0_S N_VDD_XI8.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI7.X0_PGD N_VDD_c_65_p N_VDD_c_3_p N_VDD_c_66_p N_VDD_c_6_p
+ N_VDD_c_37_p N_VDD_c_9_p N_VDD_c_31_p N_VDD_c_13_p N_VDD_c_4_p N_VDD_c_36_p
+ N_VDD_c_38_p N_VDD_c_7_p N_VDD_c_40_p N_VDD_c_11_p N_VDD_c_15_p VDD
+ N_VDD_c_33_p N_VDD_c_34_p N_VDD_c_12_p N_VDD_c_16_p Vss PM_G4_MAJ3_N1_VDD
x_PM_G4_MAJ3_N1_VSS N_VSS_XI6.X0_PGD N_VSS_XI8.X0_PGD N_VSS_XI5.X0_D
+ N_VSS_XI7.X0_S N_VSS_c_83_n N_VSS_c_85_n N_VSS_c_86_n N_VSS_c_88_n
+ N_VSS_c_135_p N_VSS_c_89_n N_VSS_c_93_n N_VSS_c_97_n N_VSS_c_98_n
+ N_VSS_c_101_n N_VSS_c_102_n N_VSS_c_106_n N_VSS_c_110_n N_VSS_c_115_n
+ N_VSS_c_117_n N_VSS_c_118_n N_VSS_c_120_n N_VSS_c_121_n N_VSS_c_122_n
+ N_VSS_c_123_n VSS Vss PM_G4_MAJ3_N1_VSS
x_PM_G4_MAJ3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI2.X0_S N_A_XI3.X0_S
+ N_A_XI3.X0_PGD N_A_XI1.X0_PGD N_A_c_182_n N_A_c_171_n N_A_c_211_p N_A_c_213_p
+ N_A_c_172_n N_A_c_189_n N_A_c_177_n N_A_c_233_p N_A_c_199_p N_A_c_237_p
+ N_A_c_225_p N_A_c_236_p N_A_c_179_n A N_A_c_180_n N_A_c_207_p Vss
+ PM_G4_MAJ3_N1_A
x_PM_G4_MAJ3_N1_BI N_BI_XI6.X0_D N_BI_XI2.X0_CG N_BI_XI1.X0_CG N_BI_c_265_n
+ N_BI_c_253_n N_BI_c_262_n N_BI_c_269_n N_BI_c_270_n N_BI_c_271_n N_BI_c_273_n
+ N_BI_c_293_p N_BI_c_296_p Vss PM_G4_MAJ3_N1_BI
x_PM_G4_MAJ3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_315_n
+ N_AI_c_316_n N_AI_c_317_n N_AI_c_320_n N_AI_c_330_n N_AI_c_321_n Vss
+ PM_G4_MAJ3_N1_AI
x_PM_G4_MAJ3_N1_B N_B_XI6.X0_CG N_B_XI5.X0_CG N_B_XI4.X0_CG N_B_XI3.X0_CG
+ N_B_c_359_n N_B_c_377_n N_B_c_414_n N_B_c_361_n B N_B_c_380_n N_B_c_381_n
+ N_B_c_364_n N_B_c_386_n N_B_c_387_n N_B_c_371_n N_B_c_372_n N_B_c_405_n
+ N_B_c_408_n N_B_c_411_n N_B_c_412_n Vss PM_G4_MAJ3_N1_B
x_PM_G4_MAJ3_N1_C N_C_XI4.X0_S N_C_XI1.X0_S N_C_c_433_n N_C_c_435_n C
+ N_C_c_437_n N_C_c_436_n Vss PM_G4_MAJ3_N1_C
x_PM_G4_MAJ3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_463_n Z Vss PM_G4_MAJ3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017247f
cc_2 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172036f
cc_3 N_VDD_c_3_p N_VSS_c_83_n 0.0017247f
cc_4 N_VDD_c_4_p N_VSS_c_83_n 2.74208e-19
cc_5 N_VDD_c_4_p N_VSS_c_85_n 3.60588e-19
cc_6 N_VDD_c_6_p N_VSS_c_86_n 0.00172036f
cc_7 N_VDD_c_7_p N_VSS_c_86_n 2.46461e-19
cc_8 N_VDD_c_7_p N_VSS_c_88_n 3.60588e-19
cc_9 N_VDD_c_9_p N_VSS_c_89_n 4.43871e-19
cc_10 N_VDD_c_4_p N_VSS_c_89_n 0.00161703f
cc_11 N_VDD_c_11_p N_VSS_c_89_n 9.28314e-19
cc_12 N_VDD_c_12_p N_VSS_c_89_n 3.48267e-19
cc_13 N_VDD_c_13_p N_VSS_c_93_n 4.43871e-19
cc_14 N_VDD_c_7_p N_VSS_c_93_n 0.00161703f
cc_15 N_VDD_c_15_p N_VSS_c_93_n 8.31866e-19
cc_16 N_VDD_c_16_p N_VSS_c_93_n 3.48267e-19
cc_17 N_VDD_c_11_p N_VSS_c_97_n 8.49247e-19
cc_18 N_VDD_XI7.X0_PGD N_VSS_c_98_n 3.41313e-19
cc_19 N_VDD_c_15_p N_VSS_c_98_n 0.00507115f
cc_20 N_VDD_c_16_p N_VSS_c_98_n 9.58524e-19
cc_21 N_VDD_c_7_p N_VSS_c_101_n 0.00403287f
cc_22 N_VDD_c_9_p N_VSS_c_102_n 3.66936e-19
cc_23 N_VDD_c_4_p N_VSS_c_102_n 2.03837e-19
cc_24 N_VDD_c_11_p N_VSS_c_102_n 3.99794e-19
cc_25 N_VDD_c_12_p N_VSS_c_102_n 8.07896e-19
cc_26 N_VDD_c_13_p N_VSS_c_106_n 3.66936e-19
cc_27 N_VDD_c_7_p N_VSS_c_106_n 2.03837e-19
cc_28 N_VDD_c_15_p N_VSS_c_106_n 3.99794e-19
cc_29 N_VDD_c_16_p N_VSS_c_106_n 8.03027e-19
cc_30 N_VDD_c_9_p N_VSS_c_110_n 0.00303537f
cc_31 N_VDD_c_31_p N_VSS_c_110_n 0.00599011f
cc_32 N_VDD_c_13_p N_VSS_c_110_n 0.00284565f
cc_33 N_VDD_c_33_p N_VSS_c_110_n 0.00104624f
cc_34 N_VDD_c_34_p N_VSS_c_110_n 0.0010706f
cc_35 N_VDD_c_4_p N_VSS_c_115_n 0.00345066f
cc_36 N_VDD_c_36_p N_VSS_c_115_n 2.07484e-19
cc_37 N_VDD_c_37_p N_VSS_c_117_n 0.00106317f
cc_38 N_VDD_c_38_p N_VSS_c_118_n 2.07484e-19
cc_39 N_VDD_c_7_p N_VSS_c_118_n 0.00345066f
cc_40 N_VDD_c_40_p N_VSS_c_120_n 0.00106317f
cc_41 N_VDD_c_4_p N_VSS_c_121_n 0.00557569f
cc_42 N_VDD_c_4_p N_VSS_c_122_n 7.74609e-19
cc_43 N_VDD_c_7_p N_VSS_c_123_n 7.74609e-19
cc_44 N_VDD_c_16_p N_A_XI7.X0_CG 9.92565e-19
cc_45 N_VDD_XI7.X0_PGD N_A_c_171_n 3.90792e-19
cc_46 N_VDD_XI7.X0_PGD N_A_c_172_n 5.17967e-19
cc_47 N_VDD_c_4_p N_A_c_172_n 3.35498e-19
cc_48 N_VDD_c_7_p N_A_c_172_n 4.32724e-19
cc_49 N_VDD_c_15_p N_A_c_172_n 4.1682e-19
cc_50 N_VDD_c_16_p N_A_c_172_n 5.53168e-19
cc_51 N_VDD_c_11_p N_A_c_177_n 5.52801e-19
cc_52 N_VDD_c_12_p N_A_c_177_n 4.1541e-19
cc_53 N_VDD_c_31_p N_A_c_179_n 5.53687e-19
cc_54 N_VDD_c_31_p N_A_c_180_n 4.71537e-19
cc_55 N_VDD_XI6.X0_S N_BI_XI6.X0_D 3.43419e-19
cc_56 N_VDD_c_4_p N_BI_XI6.X0_D 3.70842e-19
cc_57 N_VDD_c_36_p N_BI_XI6.X0_D 3.72199e-19
cc_58 N_VDD_XI6.X0_S N_BI_c_253_n 3.48267e-19
cc_59 N_VDD_c_4_p N_BI_c_253_n 4.45573e-19
cc_60 N_VDD_c_36_p N_BI_c_253_n 5.2846e-19
cc_61 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_62 N_VDD_c_38_p N_AI_XI8.X0_D 3.72199e-19
cc_63 N_VDD_XI5.X0_PGD N_AI_XI2.X0_PGD 2.73831e-19
cc_64 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.86706e-19
cc_65 N_VDD_c_65_p N_AI_c_315_n 2.73831e-19
cc_66 N_VDD_c_66_p N_AI_c_316_n 2.86706e-19
cc_67 N_VDD_XI8.X0_S N_AI_c_317_n 3.48267e-19
cc_68 N_VDD_c_38_p N_AI_c_317_n 5.226e-19
cc_69 N_VDD_c_7_p N_AI_c_317_n 5.01863e-19
cc_70 N_VDD_c_15_p N_AI_c_320_n 0.00114922f
cc_71 N_VDD_c_7_p N_AI_c_321_n 2.39469e-19
cc_72 N_VDD_c_12_p N_B_XI5.X0_CG 0.00237871f
cc_73 N_VDD_XI5.X0_PGD N_B_c_359_n 3.9688e-19
cc_74 N_VDD_XI7.X0_PGD N_B_c_359_n 2.07132e-19
cc_75 N_VDD_c_31_p N_B_c_361_n 3.8625e-19
cc_76 N_VDD_c_11_p N_B_c_361_n 6.84022e-19
cc_77 N_VDD_c_12_p N_B_c_361_n 8.63725e-19
cc_78 N_VDD_c_11_p N_B_c_364_n 4.85469e-19
cc_79 N_VDD_c_12_p N_B_c_364_n 0.0014909f
cc_80 N_VDD_c_16_p N_B_c_364_n 5.33198e-19
cc_81 N_VSS_XI5.X0_D N_A_XI2.X0_S 3.43419e-19
cc_82 N_VSS_c_106_n N_A_c_182_n 0.00236445f
cc_83 N_VSS_XI8.X0_PGD N_A_c_171_n 3.86211e-19
cc_84 N_VSS_XI7.X0_S N_A_c_172_n 9.18655e-19
cc_85 N_VSS_c_97_n N_A_c_172_n 4.08476e-19
cc_86 N_VSS_c_98_n N_A_c_172_n 0.00149476f
cc_87 N_VSS_c_101_n N_A_c_172_n 2.91598e-19
cc_88 N_VSS_c_121_n N_A_c_172_n 2.51207e-19
cc_89 N_VSS_XI5.X0_D N_A_c_189_n 9.18655e-19
cc_90 N_VSS_c_97_n N_A_c_189_n 0.00202821f
cc_91 N_VSS_c_97_n N_A_c_177_n 0.0012307f
cc_92 N_VSS_c_135_p N_A_c_179_n 3.48564e-19
cc_93 N_VSS_c_93_n N_A_c_179_n 5.0102e-19
cc_94 N_VSS_c_106_n N_A_c_179_n 4.64764e-19
cc_95 N_VSS_c_110_n N_A_c_179_n 4.46304e-19
cc_96 N_VSS_c_93_n N_A_c_180_n 4.26083e-19
cc_97 N_VSS_c_102_n N_A_c_180_n 5.39888e-19
cc_98 N_VSS_c_106_n N_A_c_180_n 0.001324f
cc_99 N_VSS_XI5.X0_D N_BI_XI6.X0_D 3.43419e-19
cc_100 N_VSS_c_97_n N_BI_XI6.X0_D 3.48267e-19
cc_101 N_VSS_XI5.X0_D N_BI_c_253_n 3.48267e-19
cc_102 N_VSS_c_97_n N_BI_c_253_n 0.0010124f
cc_103 N_VSS_c_110_n N_BI_c_253_n 6.76595e-19
cc_104 N_VSS_c_121_n N_BI_c_253_n 6.07981e-19
cc_105 N_VSS_c_97_n N_BI_c_262_n 5.26238e-19
cc_106 N_VSS_c_121_n N_BI_c_262_n 7.0632e-19
cc_107 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_108 N_VSS_c_98_n N_AI_XI8.X0_D 3.48267e-19
cc_109 N_VSS_c_98_n N_AI_XI2.X0_PGD 2.04949e-19
cc_110 N_VSS_XI7.X0_S N_AI_c_317_n 3.48267e-19
cc_111 N_VSS_c_93_n N_AI_c_317_n 0.00173262f
cc_112 N_VSS_c_98_n N_AI_c_317_n 0.00129107f
cc_113 N_VSS_c_110_n N_AI_c_317_n 9.31051e-19
cc_114 N_VSS_c_98_n N_AI_c_320_n 0.00170897f
cc_115 N_VSS_c_98_n N_AI_c_330_n 2.82216e-19
cc_116 N_VSS_c_101_n N_AI_c_321_n 0.00934196f
cc_117 N_VSS_c_102_n N_B_XI6.X0_CG 9.70552e-19
cc_118 N_VSS_XI6.X0_PGD N_B_c_359_n 3.923e-19
cc_119 N_VSS_XI8.X0_PGD N_B_c_359_n 2.07132e-19
cc_120 N_VSS_c_110_n N_B_c_361_n 7.87668e-19
cc_121 N_VSS_c_97_n N_B_c_371_n 5.49592e-19
cc_122 N_VSS_c_101_n N_B_c_372_n 2.27662e-19
cc_123 N_VSS_XI7.X0_S N_C_XI4.X0_S 3.43419e-19
cc_124 N_VSS_c_98_n N_C_XI4.X0_S 3.48267e-19
cc_125 N_VSS_XI7.X0_S N_C_c_433_n 3.48267e-19
cc_126 N_VSS_c_98_n N_C_c_433_n 5.64614e-19
cc_127 N_A_c_199_p N_BI_XI2.X0_CG 2.16788e-19
cc_128 N_A_XI3.X0_PGD N_BI_c_265_n 8.79767e-19
cc_129 N_A_c_172_n N_BI_c_253_n 0.00115944f
cc_130 N_A_c_189_n N_BI_c_262_n 0.00163472f
cc_131 N_A_c_199_p N_BI_c_262_n 0.00112713f
cc_132 N_A_c_199_p N_BI_c_269_n 5.2034e-19
cc_133 N_A_c_189_n N_BI_c_270_n 3.37713e-19
cc_134 N_A_XI3.X0_PGD N_BI_c_271_n 0.00245019f
cc_135 N_A_c_207_p N_BI_c_271_n 3.56342e-19
cc_136 N_A_c_199_p N_BI_c_273_n 0.00124805f
cc_137 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174421f
cc_138 N_A_c_189_n N_AI_XI2.X0_PGD 8.48901e-19
cc_139 N_A_c_211_p N_AI_c_315_n 0.00195894f
cc_140 N_A_c_199_p N_AI_c_315_n 0.00178666f
cc_141 N_A_c_213_p N_AI_c_316_n 0.00202303f
cc_142 N_A_c_172_n N_AI_c_317_n 0.00165136f
cc_143 N_A_c_172_n N_AI_c_320_n 0.00201403f
cc_144 N_A_XI3.X0_PGD N_B_XI3.X0_CG 8.79767e-19
cc_145 N_A_c_207_p N_B_XI3.X0_CG 0.00234701f
cc_146 N_A_c_171_n N_B_c_359_n 0.0036024f
cc_147 N_A_c_172_n N_B_c_359_n 5.44634e-19
cc_148 N_A_c_180_n N_B_c_377_n 4.18059e-19
cc_149 N_A_c_172_n N_B_c_361_n 7.76373e-19
cc_150 N_A_c_189_n N_B_c_361_n 0.00128334f
cc_151 N_A_c_172_n N_B_c_380_n 3.26436e-19
cc_152 N_A_c_199_p N_B_c_381_n 3.96409e-19
cc_153 N_A_c_225_p N_B_c_381_n 9.9319e-19
cc_154 N_A_c_207_p N_B_c_381_n 4.87397e-19
cc_155 N_A_c_171_n N_B_c_364_n 3.81736e-19
cc_156 N_A_c_189_n N_B_c_364_n 5.63683e-19
cc_157 N_A_c_172_n N_B_c_386_n 3.8563e-19
cc_158 N_A_XI3.X0_PGD N_B_c_387_n 0.00312702f
cc_159 N_A_c_207_p N_B_c_387_n 0.00145837f
cc_160 N_A_c_189_n N_B_c_371_n 0.002414f
cc_161 N_A_c_233_p N_B_c_371_n 3.98537e-19
cc_162 N_A_c_199_p N_B_c_371_n 6.08993e-19
cc_163 N_A_c_172_n N_B_c_372_n 0.00197865f
cc_164 N_A_c_236_p N_C_c_435_n 2.22411e-19
cc_165 N_A_c_237_p N_C_c_436_n 4.03103e-19
cc_166 N_A_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_167 N_A_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_168 N_A_c_233_p N_Z_XI2.X0_D 3.48267e-19
cc_169 N_A_c_199_p N_Z_XI2.X0_D 9.18655e-19
cc_170 N_A_c_236_p N_Z_XI2.X0_D 3.48267e-19
cc_171 N_A_XI2.X0_S N_Z_c_463_n 3.48267e-19
cc_172 N_A_XI3.X0_S N_Z_c_463_n 3.48267e-19
cc_173 N_A_XI3.X0_PGD N_Z_c_463_n 5.57521e-19
cc_174 N_A_c_189_n N_Z_c_463_n 9.24e-19
cc_175 N_A_c_233_p N_Z_c_463_n 7.8992e-19
cc_176 N_A_c_199_p N_Z_c_463_n 0.00158543f
cc_177 N_A_c_236_p N_Z_c_463_n 8.08848e-19
cc_178 N_BI_XI2.X0_CG N_AI_XI2.X0_PGD 8.63152e-19
cc_179 N_BI_c_270_n N_AI_XI2.X0_PGD 0.00312702f
cc_180 N_BI_c_253_n N_AI_c_317_n 3.22835e-19
cc_181 N_BI_c_262_n N_AI_c_320_n 3.68388e-19
cc_182 N_BI_c_270_n N_AI_c_330_n 2.00604e-19
cc_183 N_BI_c_262_n N_B_c_361_n 0.00136623f
cc_184 N_BI_c_262_n N_B_c_380_n 6.77523e-19
cc_185 N_BI_c_270_n N_B_c_380_n 4.99367e-19
cc_186 N_BI_c_269_n N_B_c_381_n 0.00186236f
cc_187 N_BI_c_271_n N_B_c_381_n 4.99367e-19
cc_188 N_BI_c_273_n N_B_c_381_n 0.00166575f
cc_189 N_BI_c_270_n N_B_c_386_n 0.00513784f
cc_190 N_BI_c_271_n N_B_c_386_n 7.2092e-19
cc_191 N_BI_c_269_n N_B_c_387_n 4.99367e-19
cc_192 N_BI_c_270_n N_B_c_387_n 6.22265e-19
cc_193 N_BI_c_271_n N_B_c_387_n 0.00499463f
cc_194 N_BI_c_262_n N_B_c_371_n 0.00525284f
cc_195 N_BI_c_262_n N_B_c_405_n 2.67017e-19
cc_196 N_BI_c_273_n N_B_c_405_n 0.0013533f
cc_197 N_BI_c_293_p N_B_c_405_n 0.00340518f
cc_198 N_BI_c_262_n N_B_c_408_n 4.99817e-19
cc_199 N_BI_c_273_n N_B_c_408_n 9.35879e-19
cc_200 N_BI_c_296_p N_B_c_408_n 7.59935e-19
cc_201 N_BI_c_293_p N_B_c_411_n 0.00181541f
cc_202 N_BI_c_262_n N_B_c_412_n 0.00138818f
cc_203 N_BI_c_273_n N_B_c_412_n 8.23093e-19
cc_204 N_BI_c_262_n N_C_c_437_n 3.43796e-19
cc_205 N_BI_c_262_n N_C_c_436_n 7.49861e-19
cc_206 N_BI_c_269_n N_C_c_436_n 9.95458e-19
cc_207 N_BI_c_296_p N_C_c_436_n 3.37189e-19
cc_208 N_BI_c_262_n N_Z_c_463_n 0.00187303f
cc_209 N_BI_c_269_n N_Z_c_463_n 0.00192908f
cc_210 N_BI_c_270_n N_Z_c_463_n 8.66889e-19
cc_211 N_BI_c_271_n N_Z_c_463_n 8.66889e-19
cc_212 N_BI_c_273_n N_Z_c_463_n 7.39431e-19
cc_213 N_BI_c_293_p N_Z_c_463_n 0.00210701f
cc_214 N_BI_c_296_p N_Z_c_463_n 9.92397e-19
cc_215 N_AI_XI2.X0_PGD N_B_c_414_n 8.79767e-19
cc_216 N_AI_c_330_n N_B_c_414_n 0.00234701f
cc_217 N_AI_c_320_n N_B_c_380_n 5.22873e-19
cc_218 N_AI_c_330_n N_B_c_380_n 4.87397e-19
cc_219 N_AI_XI2.X0_PGD N_B_c_386_n 0.00312702f
cc_220 N_AI_c_320_n N_B_c_386_n 4.3265e-19
cc_221 N_AI_c_330_n N_B_c_386_n 0.00145837f
cc_222 N_AI_c_320_n N_B_c_372_n 0.00441104f
cc_223 N_AI_c_320_n N_B_c_405_n 3.85994e-19
cc_224 N_AI_c_320_n N_C_c_433_n 0.00187508f
cc_225 N_AI_c_317_n N_C_c_437_n 2.87718e-19
cc_226 N_AI_c_320_n N_C_c_437_n 8.98954e-19
cc_227 N_AI_c_320_n N_C_c_436_n 5.19511e-19
cc_228 N_AI_XI2.X0_PGD N_Z_c_463_n 2.98914e-19
cc_229 N_B_c_371_n N_C_c_433_n 8.83421e-19
cc_230 N_B_c_381_n N_C_c_436_n 9.42245e-19
cc_231 N_B_c_371_n N_C_c_436_n 2.24447e-19
cc_232 N_B_c_408_n N_C_c_436_n 0.00527131f
cc_233 N_B_c_380_n N_Z_c_463_n 0.00210511f
cc_234 N_B_c_381_n N_Z_c_463_n 0.00187303f
cc_235 N_B_c_387_n N_Z_c_463_n 8.66889e-19
cc_236 N_B_c_405_n N_Z_c_463_n 4.75654e-19
cc_237 N_C_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_238 N_C_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_239 N_C_c_433_n N_Z_XI4.X0_D 3.48267e-19
cc_240 N_C_c_435_n N_Z_XI4.X0_D 3.48267e-19
cc_241 N_C_XI4.X0_S N_Z_c_463_n 3.48267e-19
cc_242 N_C_XI1.X0_S N_Z_c_463_n 3.48267e-19
cc_243 N_C_c_433_n N_Z_c_463_n 5.74266e-19
cc_244 N_C_c_435_n N_Z_c_463_n 5.79289e-19
cc_245 N_C_c_436_n N_Z_c_463_n 4.30842e-19
*
.ends
*
*
.subckt MAJ3_HPNW4 A B C Y VDD VSS
xgate (VDD VSS A B C Y) G4_MAJ3_N1_2
.ends
*
* File: G3_MIN3_T6_N1.pex.netlist
* Created: Sun Apr 10 19:28:11 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*






.subckt G3_MIN3_T6_N1_2 VSS VDD Z C B A
*
* A	A
* B	B
* C	C
* Z	Z
* VDD	VDD
* VSS	VSS
XI9.X0 N_Z_XI9.X0_D N_VSS_XI9.X0_PGD N_C_XI9.X0_CG N_B_XI9.X0_PGS N_VDD_XI9.X0_S
+ TIGFET_HPNW4
XI6.X0 N_Z_XI6.X0_D N_VDD_XI6.X0_PGD N_C_XI6.X0_CG N_B_XI6.X0_PGS N_VSS_XI6.X0_S
+ TIGFET_HPNW4
XI11.X0 N_Z_XI11.X0_D N_VSS_XI11.X0_PGD N_A_XI11.X0_CG N_B_XI11.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW4
XI10.X0 N_Z_XI10.X0_D N_VDD_XI10.X0_PGD N_A_XI10.X0_CG N_B_XI10.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW4
XI8.X0 N_Z_XI11.X0_D N_VSS_XI8.X0_PGD N_C_XI8.X0_CG N_A_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI7.X0 N_Z_XI10.X0_D N_VDD_XI7.X0_PGD N_C_XI7.X0_CG N_A_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW4
*
x_PM_G3_MIN3_T6_N1_VSS N_VSS_XI9.X0_PGD N_VSS_XI6.X0_S N_VSS_XI11.X0_PGD
+ N_VSS_XI8.X0_PGD N_VSS_XI7.X0_S N_VSS_c_8_p N_VSS_c_24_p N_VSS_c_27_p
+ N_VSS_c_9_p N_VSS_c_15_p N_VSS_c_16_p N_VSS_c_61_p N_VSS_c_10_p N_VSS_c_2_p
+ N_VSS_c_6_p N_VSS_c_11_p N_VSS_c_12_p N_VSS_c_13_p N_VSS_c_19_p N_VSS_c_28_p
+ VSS N_VSS_c_31_p N_VSS_c_76_p Vss PM_G3_MIN3_T6_N1_VSS
x_PM_G3_MIN3_T6_N1_VDD N_VDD_XI9.X0_S N_VDD_XI6.X0_PGD N_VDD_XI10.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI7.X0_PGD N_VDD_c_87_n N_VDD_c_150_p N_VDD_c_160_p
+ N_VDD_c_153_p N_VDD_c_152_p N_VDD_c_88_n N_VDD_c_93_n N_VDD_c_99_n
+ N_VDD_c_100_n N_VDD_c_102_n N_VDD_c_105_n N_VDD_c_108_n N_VDD_c_142_p VDD
+ N_VDD_c_111_n Vss PM_G3_MIN3_T6_N1_VDD
x_PM_G3_MIN3_T6_N1_Z N_Z_XI9.X0_D N_Z_XI6.X0_D N_Z_XI11.X0_D N_Z_XI10.X0_D
+ N_Z_c_170_n N_Z_c_176_n Z N_Z_c_180_n Vss PM_G3_MIN3_T6_N1_Z
x_PM_G3_MIN3_T6_N1_C N_C_XI9.X0_CG N_C_XI6.X0_CG N_C_XI8.X0_CG N_C_XI7.X0_CG
+ N_C_c_212_n N_C_c_213_n C N_C_c_214_n N_C_c_215_n N_C_c_216_n Vss
+ PM_G3_MIN3_T6_N1_C
x_PM_G3_MIN3_T6_N1_B N_B_XI9.X0_PGS N_B_XI6.X0_PGS N_B_XI11.X0_PGS
+ N_B_XI10.X0_PGS N_B_c_247_n N_B_c_248_n N_B_c_256_n B N_B_c_258_n Vss
+ PM_G3_MIN3_T6_N1_B
x_PM_G3_MIN3_T6_N1_A N_A_XI11.X0_CG N_A_XI10.X0_CG N_A_XI8.X0_PGS N_A_XI7.X0_PGS
+ N_A_c_272_n A N_A_c_276_n N_A_c_282_n N_A_c_283_n Vss PM_G3_MIN3_T6_N1_A
cc_1 N_VSS_XI6.X0_S N_VDD_XI9.X0_S 4.21365e-19
cc_2 N_VSS_c_2_p N_VDD_XI9.X0_S 3.8999e-19
cc_3 N_VSS_XI9.X0_PGD N_VDD_XI6.X0_PGD 6.1888e-19
cc_4 N_VSS_XI11.X0_PGD N_VDD_XI10.X0_PGD 6.1888e-19
cc_5 N_VSS_XI7.X0_S N_VDD_XI8.X0_S 4.21365e-19
cc_6 N_VSS_c_6_p N_VDD_XI8.X0_S 3.8999e-19
cc_7 N_VSS_XI8.X0_PGD N_VDD_XI7.X0_PGD 5.98857e-19
cc_8 N_VSS_c_8_p N_VDD_c_87_n 6.35797e-19
cc_9 N_VSS_c_9_p N_VDD_c_88_n 2.61781e-19
cc_10 N_VSS_c_10_p N_VDD_c_88_n 0.00161042f
cc_11 N_VSS_c_11_p N_VDD_c_88_n 0.00118088f
cc_12 N_VSS_c_12_p N_VDD_c_88_n 0.00296683f
cc_13 N_VSS_c_13_p N_VDD_c_88_n 0.00183744f
cc_14 N_VSS_c_9_p N_VDD_c_93_n 9.27292e-19
cc_15 N_VSS_c_15_p N_VDD_c_93_n 3.72495e-19
cc_16 N_VSS_c_16_p N_VDD_c_93_n 8.87931e-19
cc_17 N_VSS_c_10_p N_VDD_c_93_n 9.0356e-19
cc_18 N_VSS_c_11_p N_VDD_c_93_n 4.3265e-19
cc_19 N_VSS_c_19_p N_VDD_c_93_n 3.0156e-19
cc_20 N_VSS_c_12_p N_VDD_c_99_n 0.00167687f
cc_21 N_VSS_c_10_p N_VDD_c_100_n 0.00121886f
cc_22 N_VSS_c_19_p N_VDD_c_100_n 3.71304e-19
cc_23 N_VSS_XI6.X0_S N_VDD_c_102_n 4.24828e-19
cc_24 N_VSS_c_24_p N_VDD_c_102_n 0.00115189f
cc_25 N_VSS_c_2_p N_VDD_c_102_n 4.59126e-19
cc_26 N_VSS_c_24_p N_VDD_c_105_n 9.72233e-19
cc_27 N_VSS_c_27_p N_VDD_c_105_n 8.14547e-19
cc_28 N_VSS_c_28_p N_VDD_c_105_n 3.32851e-19
cc_29 N_VSS_XI7.X0_S N_VDD_c_108_n 3.8999e-19
cc_30 N_VSS_c_6_p N_VDD_c_108_n 5.78716e-19
cc_31 N_VSS_c_31_p N_VDD_c_108_n 0.00180659f
cc_32 N_VSS_c_10_p N_VDD_c_111_n 3.8999e-19
cc_33 N_VSS_c_11_p N_VDD_c_111_n 0.00181085f
cc_34 N_VSS_c_10_p N_Z_XI9.X0_D 8.835e-19
cc_35 N_VSS_c_11_p N_Z_XI9.X0_D 0.00246958f
cc_36 N_VSS_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_37 N_VSS_c_2_p N_Z_XI6.X0_D 3.48267e-19
cc_38 N_VSS_XI6.X0_S N_Z_XI10.X0_D 3.43419e-19
cc_39 N_VSS_XI7.X0_S N_Z_XI10.X0_D 3.43419e-19
cc_40 N_VSS_c_2_p N_Z_XI10.X0_D 3.48267e-19
cc_41 N_VSS_c_6_p N_Z_XI10.X0_D 3.48267e-19
cc_42 N_VSS_XI6.X0_S N_Z_c_170_n 3.48267e-19
cc_43 N_VSS_c_10_p N_Z_c_170_n 0.00217565f
cc_44 N_VSS_c_2_p N_Z_c_170_n 5.69026e-19
cc_45 N_VSS_c_11_p N_Z_c_170_n 8.835e-19
cc_46 N_VSS_c_12_p N_Z_c_170_n 7.10715e-19
cc_47 N_VSS_c_19_p N_Z_c_170_n 3.30259e-19
cc_48 N_VSS_XI6.X0_S N_Z_c_176_n 3.48267e-19
cc_49 N_VSS_XI7.X0_S N_Z_c_176_n 3.48267e-19
cc_50 N_VSS_c_2_p N_Z_c_176_n 5.69026e-19
cc_51 N_VSS_c_6_p N_Z_c_176_n 5.69026e-19
cc_52 N_VSS_c_2_p N_Z_c_180_n 0.00191849f
cc_53 N_VSS_c_12_p N_Z_c_180_n 5.57576e-19
cc_54 N_VSS_c_19_p N_Z_c_180_n 0.00201399f
cc_55 N_VSS_c_28_p N_Z_c_180_n 5.26184e-19
cc_56 N_VSS_XI9.X0_PGD N_C_c_212_n 4.30517e-19
cc_57 N_VSS_XI8.X0_PGD N_C_c_213_n 5.02359e-19
cc_58 N_VSS_c_28_p N_C_c_214_n 2.73385e-19
cc_59 N_VSS_XI9.X0_PGD N_C_c_215_n 4.3583e-19
cc_60 N_VSS_XI8.X0_PGD N_C_c_216_n 3.76133e-19
cc_61 N_VSS_c_61_p N_C_c_216_n 2.17009e-19
cc_62 N_VSS_XI9.X0_PGD N_B_XI9.X0_PGS 0.00109504f
cc_63 N_VSS_XI11.X0_PGD N_B_XI9.X0_PGS 2.15671e-19
cc_64 N_VSS_XI11.X0_PGD N_B_XI11.X0_PGS 0.00177732f
cc_65 N_VSS_XI8.X0_PGD N_B_XI11.X0_PGS 2.22194e-19
cc_66 N_VSS_c_61_p N_B_c_247_n 0.00177732f
cc_67 N_VSS_c_24_p N_B_c_248_n 0.00731987f
cc_68 N_VSS_c_16_p N_B_c_248_n 0.00109504f
cc_69 N_VSS_c_2_p B 2.11465e-19
cc_70 N_VSS_c_12_p B 2.74582e-19
cc_71 N_VSS_c_19_p B 2.99651e-19
cc_72 N_VSS_c_24_p N_A_XI11.X0_CG 2.66861e-19
cc_73 N_VSS_c_2_p N_A_c_272_n 3.13396e-19
cc_74 N_VSS_c_28_p N_A_c_272_n 5.88825e-19
cc_75 N_VSS_c_28_p A 5.88825e-19
cc_76 N_VSS_c_76_p A 2.39495e-19
cc_77 N_VSS_c_2_p N_A_c_276_n 0.00159849f
cc_78 N_VSS_c_28_p N_A_c_276_n 0.00924443f
cc_79 N_VSS_c_76_p N_A_c_276_n 5.12768e-19
cc_80 N_VDD_XI9.X0_S N_Z_XI9.X0_D 3.43419e-19
cc_81 N_VDD_c_93_n N_Z_XI9.X0_D 4.3265e-19
cc_82 N_VDD_c_102_n N_Z_XI9.X0_D 3.48267e-19
cc_83 N_VDD_c_100_n N_Z_XI6.X0_D 9.44213e-19
cc_84 N_VDD_c_111_n N_Z_XI6.X0_D 0.00246958f
cc_85 N_VDD_XI9.X0_S N_Z_XI11.X0_D 3.43419e-19
cc_86 N_VDD_XI8.X0_S N_Z_XI11.X0_D 3.43419e-19
cc_87 N_VDD_c_102_n N_Z_XI11.X0_D 3.48267e-19
cc_88 N_VDD_c_105_n N_Z_XI11.X0_D 4.3265e-19
cc_89 N_VDD_c_108_n N_Z_XI11.X0_D 3.72199e-19
cc_90 N_VDD_XI9.X0_S N_Z_c_170_n 3.48267e-19
cc_91 N_VDD_c_88_n N_Z_c_170_n 0.0013145f
cc_92 N_VDD_c_93_n N_Z_c_170_n 7.37531e-19
cc_93 N_VDD_c_100_n N_Z_c_170_n 0.00186578f
cc_94 N_VDD_c_102_n N_Z_c_170_n 7.73813e-19
cc_95 N_VDD_c_111_n N_Z_c_170_n 8.835e-19
cc_96 N_VDD_XI9.X0_S N_Z_c_176_n 3.48267e-19
cc_97 N_VDD_XI8.X0_S N_Z_c_176_n 3.48267e-19
cc_98 N_VDD_c_102_n N_Z_c_176_n 8.00908e-19
cc_99 N_VDD_c_105_n N_Z_c_176_n 5.78499e-19
cc_100 N_VDD_c_108_n N_Z_c_176_n 8.53368e-19
cc_101 N_VDD_c_93_n N_Z_c_180_n 8.36802e-19
cc_102 N_VDD_c_88_n C 2.63478e-19
cc_103 N_VDD_c_93_n C 0.00145322f
cc_104 N_VDD_c_102_n C 0.00155931f
cc_105 N_VDD_c_88_n N_C_c_214_n 2.14517e-19
cc_106 N_VDD_c_93_n N_C_c_214_n 8.61717e-19
cc_107 N_VDD_c_102_n N_C_c_214_n 0.00183615f
cc_108 N_VDD_c_105_n N_C_c_214_n 0.00557625f
cc_109 N_VDD_c_142_p N_C_c_214_n 5.42852e-19
cc_110 N_VDD_c_93_n N_C_c_215_n 7.51813e-19
cc_111 N_VDD_c_102_n N_C_c_215_n 8.66889e-19
cc_112 N_VDD_c_102_n N_C_c_216_n 2.22969e-19
cc_113 N_VDD_c_105_n N_C_c_216_n 2.63125e-19
cc_114 N_VDD_c_142_p N_C_c_216_n 3.66936e-19
cc_115 N_VDD_XI6.X0_PGD N_B_XI9.X0_PGS 0.00135245f
cc_116 N_VDD_XI10.X0_PGD N_B_XI9.X0_PGS 4.12959e-19
cc_117 N_VDD_c_150_p N_B_XI11.X0_PGS 0.00109105f
cc_118 N_VDD_c_150_p N_B_c_256_n 0.00258419f
cc_119 N_VDD_c_152_p N_B_c_256_n 4.12959e-19
cc_120 N_VDD_c_153_p N_B_c_258_n 0.00495207f
cc_121 N_VDD_c_111_n N_B_c_258_n 4.60491e-19
cc_122 N_VDD_XI10.X0_PGD N_A_XI11.X0_CG 4.83278e-19
cc_123 N_VDD_XI7.X0_PGD N_A_XI8.X0_PGS 0.00141985f
cc_124 N_VDD_c_105_n N_A_XI8.X0_PGS 2.26738e-19
cc_125 N_VDD_XI10.X0_PGD N_A_c_282_n 5.50272e-19
cc_126 N_VDD_XI7.X0_PGD N_A_c_283_n 3.23173e-19
cc_127 N_VDD_c_160_p N_A_c_283_n 0.00145458f
cc_128 N_VDD_c_152_p N_A_c_283_n 2.17009e-19
cc_129 N_Z_c_170_n N_C_c_212_n 6.18749e-19
cc_130 N_Z_c_176_n N_C_c_213_n 8.38264e-19
cc_131 N_Z_c_180_n N_C_c_214_n 0.0071108f
cc_132 N_Z_c_176_n N_A_XI11.X0_CG 2.49716e-19
cc_133 N_Z_c_176_n N_A_c_276_n 3.55289e-19
cc_134 N_Z_c_180_n N_A_c_276_n 0.00276659f
cc_135 N_C_c_212_n N_B_XI9.X0_PGS 0.00830899f
cc_136 N_C_c_215_n N_B_XI9.X0_PGS 3.76133e-19
cc_137 N_C_c_212_n N_B_XI11.X0_PGS 8.90713e-19
cc_138 N_C_c_213_n N_B_XI11.X0_PGS 5.42381e-19
cc_139 N_C_c_215_n N_B_c_258_n 3.15193e-19
cc_140 N_C_c_213_n N_A_XI11.X0_CG 0.0020589f
cc_141 N_C_c_213_n N_A_XI8.X0_PGS 0.00810452f
cc_142 N_C_c_214_n N_A_c_276_n 0.00121525f
cc_143 N_C_c_216_n N_A_c_283_n 3.16599e-19
cc_144 N_B_XI9.X0_PGS N_A_XI11.X0_CG 0.00106357f
cc_145 N_B_XI11.X0_PGS N_A_XI11.X0_CG 0.00765248f
cc_146 B N_A_c_272_n 3.39698e-19
cc_147 N_B_c_258_n N_A_c_272_n 3.48267e-19
cc_148 B N_A_c_282_n 3.48267e-19
cc_149 N_B_c_258_n N_A_c_282_n 5.15124e-19
*
.ends
*
*
.subckt MIN3_HPNW4 A B C Y VDD VSS
xgate (VSS VDD Y C B A) G3_MIN3_T6_N1_2
.ends
*
* File: G4_MUX2_N1.pex.netlist
* Created: Wed Mar  9 17:10:36 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*








.subckt G4_MUX2_N1_2 VDD VSS Z SEL B A
*
* A	A
* B	B
* SEL	SEL
* Z	Z
* VSS	VSS
* VDD	VDD
XI7.X0 N_VDD_XI7.X0_D N_VSS_XI7.X0_PGD N_ZI_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_Z_XI7.X0_S TIGFET_HPNW4
XI1.X0 N_SELI_XI1.X0_D N_VDD_XI1.X0_PGD N_SEL_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI6.X0 N_Z_XI7.X0_S N_VDD_XI6.X0_PGD N_ZI_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW4
XI2.X0 N_SELI_XI1.X0_D N_VSS_XI2.X0_PGD N_SEL_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI5.X0 N_ZI_XI5.X0_D N_VDD_XI5.X0_PGD N_SELI_XI5.X0_CG N_B_XI5.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW4
XI3.X0 N_ZI_XI3.X0_D N_VSS_XI3.X0_PGD N_SEL_XI3.X0_CG N_B_XI3.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI4.X0 N_ZI_XI5.X0_D N_VDD_XI4.X0_PGD N_SEL_XI4.X0_CG N_A_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW4
XI0.X0 N_ZI_XI3.X0_D N_VSS_XI0.X0_PGD N_SELI_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW4
*
x_PM_G4_MUX2_N1_VDD N_VDD_XI7.X0_D N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS
+ N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI2.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_14_p N_VDD_c_11_p N_VDD_c_136_p
+ N_VDD_c_18_p N_VDD_c_12_p N_VDD_c_46_p N_VDD_c_17_p N_VDD_c_22_p N_VDD_c_15_p
+ N_VDD_c_48_p N_VDD_c_20_p N_VDD_c_3_p N_VDD_c_6_p N_VDD_c_16_p N_VDD_c_28_p
+ N_VDD_c_8_p N_VDD_c_34_p N_VDD_c_9_p N_VDD_c_32_p VDD N_VDD_c_51_p
+ N_VDD_c_55_p N_VDD_c_58_p N_VDD_c_65_p N_VDD_c_25_p N_VDD_c_21_p N_VDD_c_95_p
+ Vss PM_G4_MUX2_N1_VDD
x_PM_G4_MUX2_N1_VSS N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS N_VSS_XI1.X0_S
+ N_VSS_XI6.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS N_VSS_XI3.X0_PGD
+ N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_151_n N_VSS_c_153_n N_VSS_c_265_p
+ N_VSS_c_154_n N_VSS_c_257_p N_VSS_c_156_n N_VSS_c_157_n N_VSS_c_158_n
+ N_VSS_c_162_n N_VSS_c_166_n N_VSS_c_170_n N_VSS_c_173_n N_VSS_c_176_n
+ N_VSS_c_180_n N_VSS_c_184_n N_VSS_c_185_n N_VSS_c_186_n N_VSS_c_187_n
+ N_VSS_c_189_n N_VSS_c_192_n N_VSS_c_193_n N_VSS_c_196_n N_VSS_c_199_n
+ N_VSS_c_200_n N_VSS_c_201_n N_VSS_c_202_n VSS N_VSS_c_206_n N_VSS_c_207_n
+ N_VSS_c_208_n N_VSS_c_209_n Vss PM_G4_MUX2_N1_VSS
x_PM_G4_MUX2_N1_ZI N_ZI_XI7.X0_CG N_ZI_XI6.X0_CG N_ZI_XI5.X0_D N_ZI_XI3.X0_D
+ N_ZI_c_278_n N_ZI_c_294_n N_ZI_c_280_n N_ZI_c_282_n N_ZI_c_287_n N_ZI_c_288_n
+ N_ZI_c_311_n N_ZI_c_326_p Vss PM_G4_MUX2_N1_ZI
x_PM_G4_MUX2_N1_Z N_Z_XI7.X0_S Z Vss PM_G4_MUX2_N1_Z
x_PM_G4_MUX2_N1_SELI N_SELI_XI1.X0_D N_SELI_XI5.X0_CG N_SELI_XI0.X0_CG
+ N_SELI_c_371_n N_SELI_c_356_n N_SELI_c_359_n N_SELI_c_387_n N_SELI_c_364_n
+ N_SELI_c_365_n N_SELI_c_367_n N_SELI_c_379_n N_SELI_c_381_n N_SELI_c_395_n
+ N_SELI_c_398_n Vss PM_G4_MUX2_N1_SELI
x_PM_G4_MUX2_N1_SEL N_SEL_XI1.X0_CG N_SEL_XI2.X0_CG N_SEL_XI3.X0_CG
+ N_SEL_XI4.X0_CG N_SEL_c_434_n N_SEL_c_460_n N_SEL_c_449_n N_SEL_c_495_p
+ N_SEL_c_436_n SEL N_SEL_c_438_n N_SEL_c_439_n N_SEL_c_440_n N_SEL_c_465_n
+ N_SEL_c_453_n N_SEL_c_468_n N_SEL_c_442_n N_SEL_c_443_n N_SEL_c_444_n
+ N_SEL_c_445_n Vss PM_G4_MUX2_N1_SEL
x_PM_G4_MUX2_N1_B N_B_XI5.X0_PGS N_B_XI3.X0_PGS N_B_c_518_n B N_B_c_514_n Vss
+ PM_G4_MUX2_N1_B
x_PM_G4_MUX2_N1_A N_A_XI4.X0_PGS N_A_XI0.X0_PGS N_A_c_544_n A N_A_c_550_n Vss
+ PM_G4_MUX2_N1_A
cc_1 N_VDD_XI1.X0_PGS N_VSS_XI7.X0_PGD 2.27468e-19
cc_2 N_VDD_XI6.X0_PGD N_VSS_XI7.X0_PGS 0.00173038f
cc_3 N_VDD_c_3_p N_VSS_XI6.X0_S 3.7884e-19
cc_4 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.0016786f
cc_5 N_VDD_XI6.X0_PGS N_VSS_XI2.X0_PGS 2.11937e-19
cc_6 N_VDD_c_6_p N_VSS_XI2.X0_PGS 2.56778e-19
cc_7 N_VDD_XI5.X0_PGD N_VSS_XI3.X0_PGD 2.1536e-19
cc_8 N_VDD_c_8_p N_VSS_XI4.X0_S 3.7884e-19
cc_9 N_VDD_c_9_p N_VSS_XI4.X0_S 9.5668e-19
cc_10 N_VDD_XI4.X0_PGD N_VSS_XI0.X0_PGD 2.1536e-19
cc_11 N_VDD_c_11_p N_VSS_c_151_n 0.00173038f
cc_12 N_VDD_c_12_p N_VSS_c_151_n 3.60588e-19
cc_13 N_VDD_c_12_p N_VSS_c_153_n 3.80388e-19
cc_14 N_VDD_c_14_p N_VSS_c_154_n 0.0016786f
cc_15 N_VDD_c_15_p N_VSS_c_154_n 2.72324e-19
cc_16 N_VDD_c_16_p N_VSS_c_156_n 8.01165e-19
cc_17 N_VDD_c_17_p N_VSS_c_157_n 9.30123e-19
cc_18 N_VDD_c_18_p N_VSS_c_158_n 8.69498e-19
cc_19 N_VDD_c_12_p N_VSS_c_158_n 0.00141228f
cc_20 N_VDD_c_20_p N_VSS_c_158_n 8.51944e-19
cc_21 N_VDD_c_21_p N_VSS_c_158_n 3.48267e-19
cc_22 N_VDD_c_22_p N_VSS_c_162_n 8.56577e-19
cc_23 N_VDD_c_15_p N_VSS_c_162_n 0.00141228f
cc_24 N_VDD_c_6_p N_VSS_c_162_n 0.00181129f
cc_25 N_VDD_c_25_p N_VSS_c_162_n 3.48267e-19
cc_26 N_VDD_c_20_p N_VSS_c_166_n 3.92901e-19
cc_27 N_VDD_c_3_p N_VSS_c_166_n 4.58491e-19
cc_28 N_VDD_c_28_p N_VSS_c_166_n 7.06793e-19
cc_29 N_VDD_c_9_p N_VSS_c_166_n 2.71563e-19
cc_30 N_VDD_c_6_p N_VSS_c_170_n 2.93442e-19
cc_31 N_VDD_c_16_p N_VSS_c_170_n 0.00161703f
cc_32 N_VDD_c_32_p N_VSS_c_170_n 4.6996e-19
cc_33 N_VDD_c_8_p N_VSS_c_173_n 4.73473e-19
cc_34 N_VDD_c_34_p N_VSS_c_173_n 2.13058e-19
cc_35 N_VDD_c_9_p N_VSS_c_173_n 0.00165395f
cc_36 N_VDD_c_18_p N_VSS_c_176_n 3.66936e-19
cc_37 N_VDD_c_12_p N_VSS_c_176_n 0.00112249f
cc_38 N_VDD_c_20_p N_VSS_c_176_n 3.99794e-19
cc_39 N_VDD_c_21_p N_VSS_c_176_n 8.07896e-19
cc_40 N_VDD_c_22_p N_VSS_c_180_n 3.82294e-19
cc_41 N_VDD_c_15_p N_VSS_c_180_n 0.00112249f
cc_42 N_VDD_c_6_p N_VSS_c_180_n 9.55349e-19
cc_43 N_VDD_c_25_p N_VSS_c_180_n 8.0279e-19
cc_44 N_VDD_c_16_p N_VSS_c_184_n 2.03837e-19
cc_45 N_VDD_c_22_p N_VSS_c_185_n 3.85245e-19
cc_46 N_VDD_c_46_p N_VSS_c_186_n 4.93614e-19
cc_47 N_VDD_c_15_p N_VSS_c_187_n 0.003995f
cc_48 N_VDD_c_48_p N_VSS_c_187_n 0.00163298f
cc_49 N_VDD_c_12_p N_VSS_c_189_n 0.00401122f
cc_50 N_VDD_c_3_p N_VSS_c_189_n 0.0013091f
cc_51 N_VDD_c_51_p N_VSS_c_189_n 0.0010079f
cc_52 N_VDD_c_12_p N_VSS_c_192_n 0.00176255f
cc_53 N_VDD_c_15_p N_VSS_c_193_n 0.00131941f
cc_54 N_VDD_c_16_p N_VSS_c_193_n 0.00593836f
cc_55 N_VDD_c_55_p N_VSS_c_193_n 0.00111239f
cc_56 N_VDD_c_3_p N_VSS_c_196_n 0.0013091f
cc_57 N_VDD_c_8_p N_VSS_c_196_n 0.00841532f
cc_58 N_VDD_c_58_p N_VSS_c_196_n 9.6871e-19
cc_59 N_VDD_c_16_p N_VSS_c_199_n 0.00454933f
cc_60 N_VDD_c_34_p N_VSS_c_200_n 5.34009e-19
cc_61 N_VDD_c_9_p N_VSS_c_201_n 0.00304617f
cc_62 N_VDD_c_6_p N_VSS_c_202_n 2.5062e-19
cc_63 N_VDD_c_9_p N_VSS_c_202_n 0.00529507f
cc_64 N_VDD_c_32_p N_VSS_c_202_n 0.00267625f
cc_65 N_VDD_c_65_p N_VSS_c_202_n 0.0010706f
cc_66 N_VDD_c_15_p N_VSS_c_206_n 7.74609e-19
cc_67 N_VDD_c_3_p N_VSS_c_207_n 0.00104966f
cc_68 N_VDD_c_16_p N_VSS_c_208_n 7.61747e-19
cc_69 N_VDD_c_9_p N_VSS_c_209_n 8.91588e-19
cc_70 N_VDD_c_21_p N_ZI_XI6.X0_CG 9.92565e-19
cc_71 N_VDD_XI2.X0_S N_ZI_XI3.X0_D 3.43419e-19
cc_72 N_VDD_XI0.X0_S N_ZI_XI3.X0_D 3.43419e-19
cc_73 N_VDD_c_6_p N_ZI_XI3.X0_D 3.48267e-19
cc_74 N_VDD_c_34_p N_ZI_XI3.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_PGD N_ZI_c_278_n 2.22031e-19
cc_76 N_VDD_XI6.X0_PGD N_ZI_c_278_n 3.91104e-19
cc_77 N_VDD_c_8_p N_ZI_c_280_n 5.01863e-19
cc_78 N_VDD_c_9_p N_ZI_c_280_n 4.66891e-19
cc_79 N_VDD_XI2.X0_S N_ZI_c_282_n 3.48267e-19
cc_80 N_VDD_XI0.X0_S N_ZI_c_282_n 3.48267e-19
cc_81 N_VDD_c_6_p N_ZI_c_282_n 4.97272e-19
cc_82 N_VDD_c_16_p N_ZI_c_282_n 5.01863e-19
cc_83 N_VDD_c_34_p N_ZI_c_282_n 5.226e-19
cc_84 N_VDD_c_25_p N_ZI_c_287_n 5.3845e-19
cc_85 N_VDD_c_15_p N_ZI_c_288_n 3.65425e-19
cc_86 N_VDD_XI7.X0_D N_Z_XI7.X0_S 3.43419e-19
cc_87 N_VDD_c_12_p N_Z_XI7.X0_S 3.7884e-19
cc_88 N_VDD_c_17_p N_Z_XI7.X0_S 3.72199e-19
cc_89 N_VDD_XI7.X0_D Z 3.48267e-19
cc_90 N_VDD_c_12_p Z 5.12447e-19
cc_91 N_VDD_c_17_p Z 7.4527e-19
cc_92 N_VDD_XI2.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_93 N_VDD_c_15_p N_SELI_XI1.X0_D 3.7884e-19
cc_94 N_VDD_c_6_p N_SELI_XI1.X0_D 3.48267e-19
cc_95 N_VDD_c_95_p N_SELI_XI5.X0_CG 0.00237871f
cc_96 N_VDD_XI2.X0_S N_SELI_c_356_n 3.48267e-19
cc_97 N_VDD_c_15_p N_SELI_c_356_n 5.34458e-19
cc_98 N_VDD_c_6_p N_SELI_c_356_n 6.883e-19
cc_99 N_VDD_XI6.X0_PGD N_SELI_c_359_n 2.27908e-19
cc_100 N_VDD_c_15_p N_SELI_c_359_n 2.61043e-19
cc_101 N_VDD_c_20_p N_SELI_c_359_n 5.3241e-19
cc_102 N_VDD_c_3_p N_SELI_c_359_n 2.36369e-19
cc_103 N_VDD_c_21_p N_SELI_c_359_n 3.99122e-19
cc_104 N_VDD_c_9_p N_SELI_c_364_n 4.30008e-19
cc_105 N_VDD_c_28_p N_SELI_c_365_n 7.54639e-19
cc_106 N_VDD_c_95_p N_SELI_c_365_n 5.0614e-19
cc_107 N_VDD_c_28_p N_SELI_c_367_n 4.85469e-19
cc_108 N_VDD_c_95_p N_SELI_c_367_n 0.0014909f
cc_109 N_VDD_c_25_p N_SEL_XI1.X0_CG 9.92565e-19
cc_110 N_VDD_XI1.X0_PGD N_SEL_c_434_n 4.04053e-19
cc_111 N_VDD_XI6.X0_PGD N_SEL_c_434_n 2.07349e-19
cc_112 N_VDD_XI2.X0_S N_SEL_c_436_n 9.18655e-19
cc_113 N_VDD_c_6_p N_SEL_c_436_n 0.00151457f
cc_114 N_VDD_c_16_p N_SEL_c_438_n 4.35337e-19
cc_115 N_VDD_c_9_p N_SEL_c_439_n 4.25334e-19
cc_116 N_VDD_c_16_p N_SEL_c_440_n 2.49768e-19
cc_117 N_VDD_c_8_p N_SEL_c_440_n 4.35337e-19
cc_118 N_VDD_c_9_p N_SEL_c_442_n 8.17234e-19
cc_119 N_VDD_c_21_p N_SEL_c_443_n 4.93609e-19
cc_120 N_VDD_c_95_p N_SEL_c_444_n 2.00604e-19
cc_121 N_VDD_XI4.X0_PGD N_SEL_c_445_n 3.11814e-19
cc_122 N_VDD_c_9_p N_SEL_c_445_n 3.66936e-19
cc_123 N_VDD_c_6_p N_B_XI5.X0_PGS 2.48132e-19
cc_124 N_VDD_c_6_p B 0.0014278f
cc_125 N_VDD_c_16_p B 0.00141439f
cc_126 N_VDD_c_6_p N_B_c_514_n 9.67317e-19
cc_127 N_VDD_c_16_p N_B_c_514_n 0.00117371f
cc_128 N_VDD_XI4.X0_PGD N_A_XI4.X0_PGS 0.00162178f
cc_129 N_VDD_c_9_p N_A_XI4.X0_PGS 9.35727e-19
cc_130 N_VDD_c_8_p N_A_c_544_n 3.3974e-19
cc_131 N_VDD_c_9_p N_A_c_544_n 4.15738e-19
cc_132 N_VDD_c_28_p A 5.43314e-19
cc_133 N_VDD_c_8_p A 0.00141439f
cc_134 N_VDD_c_9_p A 5.30212e-19
cc_135 N_VDD_c_95_p A 3.48267e-19
cc_136 N_VDD_c_136_p N_A_c_550_n 0.00480616f
cc_137 N_VDD_c_28_p N_A_c_550_n 4.04186e-19
cc_138 N_VDD_c_8_p N_A_c_550_n 0.00117371f
cc_139 N_VDD_c_9_p N_A_c_550_n 3.66936e-19
cc_140 N_VDD_c_95_p N_A_c_550_n 6.39485e-19
cc_141 N_VSS_c_176_n N_ZI_XI7.X0_CG 0.00234241f
cc_142 N_VSS_XI6.X0_S N_ZI_XI5.X0_D 3.43419e-19
cc_143 N_VSS_XI4.X0_S N_ZI_XI5.X0_D 3.43419e-19
cc_144 N_VSS_c_173_n N_ZI_XI5.X0_D 3.48267e-19
cc_145 N_VSS_XI7.X0_PGS N_ZI_c_278_n 3.99472e-19
cc_146 N_VSS_c_158_n N_ZI_c_294_n 0.00126951f
cc_147 N_VSS_c_176_n N_ZI_c_294_n 8.72558e-19
cc_148 N_VSS_XI6.X0_S N_ZI_c_280_n 3.48267e-19
cc_149 N_VSS_XI4.X0_S N_ZI_c_280_n 3.48267e-19
cc_150 N_VSS_c_166_n N_ZI_c_280_n 0.00100597f
cc_151 N_VSS_c_173_n N_ZI_c_280_n 4.40384e-19
cc_152 N_VSS_c_196_n N_ZI_c_280_n 5.12922e-19
cc_153 N_VSS_c_200_n N_ZI_c_280_n 6.1924e-19
cc_154 N_VSS_c_202_n N_ZI_c_280_n 0.00113121f
cc_155 N_VSS_c_193_n N_ZI_c_282_n 5.12922e-19
cc_156 N_VSS_c_158_n N_ZI_c_287_n 4.56568e-19
cc_157 N_VSS_c_176_n N_ZI_c_287_n 0.0014909f
cc_158 N_VSS_c_162_n N_ZI_c_288_n 4.17431e-19
cc_159 N_VSS_c_166_n N_ZI_c_288_n 6.40656e-19
cc_160 N_VSS_c_189_n N_ZI_c_288_n 0.00101727f
cc_161 N_VSS_c_193_n N_ZI_c_288_n 0.00147997f
cc_162 N_VSS_c_196_n N_ZI_c_288_n 2.59546e-19
cc_163 N_VSS_c_187_n N_ZI_c_311_n 0.0011789f
cc_164 N_VSS_XI6.X0_S N_Z_XI7.X0_S 3.43419e-19
cc_165 N_VSS_c_166_n N_Z_XI7.X0_S 3.48267e-19
cc_166 N_VSS_XI6.X0_S Z 3.48267e-19
cc_167 N_VSS_c_166_n Z 7.85754e-19
cc_168 N_VSS_XI1.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_169 N_VSS_c_157_n N_SELI_XI1.X0_D 3.48267e-19
cc_170 N_VSS_c_184_n N_SELI_c_371_n 0.00234241f
cc_171 N_VSS_c_157_n N_SELI_c_356_n 6.0686e-19
cc_172 N_VSS_c_166_n N_SELI_c_359_n 0.00130595f
cc_173 N_VSS_c_189_n N_SELI_c_359_n 4.10258e-19
cc_174 N_VSS_c_170_n N_SELI_c_364_n 0.00135778f
cc_175 N_VSS_c_184_n N_SELI_c_364_n 4.99367e-19
cc_176 N_VSS_c_196_n N_SELI_c_364_n 4.69529e-19
cc_177 N_VSS_c_202_n N_SELI_c_364_n 9.62347e-19
cc_178 N_VSS_c_170_n N_SELI_c_379_n 4.56568e-19
cc_179 N_VSS_c_184_n N_SELI_c_379_n 0.0014909f
cc_180 N_VSS_c_196_n N_SELI_c_381_n 7.6099e-19
cc_181 N_VSS_c_202_n N_SELI_c_381_n 6.2582e-19
cc_182 N_VSS_XI7.X0_PGS N_SEL_c_434_n 2.22031e-19
cc_183 N_VSS_XI2.X0_PGD N_SEL_c_434_n 3.91879e-19
cc_184 N_VSS_c_180_n N_SEL_c_449_n 0.00272336f
cc_185 N_VSS_c_193_n N_SEL_c_436_n 4.08267e-19
cc_186 N_VSS_c_202_n N_SEL_c_439_n 2.03139e-19
cc_187 N_VSS_c_196_n N_SEL_c_440_n 2.53418e-19
cc_188 N_VSS_c_257_p N_SEL_c_453_n 3.73191e-19
cc_189 N_VSS_c_162_n N_SEL_c_453_n 6.21258e-19
cc_190 N_VSS_c_162_n N_SEL_c_443_n 4.56568e-19
cc_191 N_VSS_c_180_n N_SEL_c_443_n 0.0014909f
cc_192 N_VSS_XI3.X0_PGD N_SEL_c_444_n 3.11814e-19
cc_193 N_VSS_c_184_n N_SEL_c_445_n 2.00604e-19
cc_194 N_VSS_XI2.X0_PGS N_B_XI5.X0_PGS 0.00172969f
cc_195 N_VSS_XI3.X0_PGD N_B_XI5.X0_PGS 0.00152606f
cc_196 N_VSS_c_265_p N_B_c_518_n 0.00172969f
cc_197 N_VSS_c_170_n B 3.98896e-19
cc_198 N_VSS_c_184_n B 3.5189e-19
cc_199 N_VSS_c_156_n N_B_c_514_n 0.00295829f
cc_200 N_VSS_c_170_n N_B_c_514_n 3.5189e-19
cc_201 N_VSS_c_180_n N_B_c_514_n 7.89771e-19
cc_202 N_VSS_c_184_n N_B_c_514_n 6.80896e-19
cc_203 N_VSS_c_196_n A 2.11858e-19
cc_204 N_ZI_c_282_n N_SELI_c_356_n 3.26181e-19
cc_205 N_ZI_c_288_n N_SELI_c_356_n 0.00213954f
cc_206 N_ZI_c_278_n N_SELI_c_359_n 4.92356e-19
cc_207 N_ZI_c_288_n N_SELI_c_359_n 0.00182433f
cc_208 N_ZI_c_278_n N_SELI_c_387_n 2.38253e-19
cc_209 N_ZI_c_294_n N_SELI_c_387_n 0.00150231f
cc_210 N_ZI_c_287_n N_SELI_c_387_n 0.00110082f
cc_211 N_ZI_c_282_n N_SELI_c_364_n 0.00173524f
cc_212 N_ZI_c_280_n N_SELI_c_365_n 0.00183505f
cc_213 N_ZI_c_288_n N_SELI_c_365_n 0.00144518f
cc_214 N_ZI_c_280_n N_SELI_c_381_n 7.38292e-19
cc_215 N_ZI_c_288_n N_SELI_c_381_n 7.7914e-19
cc_216 N_ZI_c_280_n N_SELI_c_395_n 5.82645e-19
cc_217 N_ZI_c_282_n N_SELI_c_395_n 3.22755e-19
cc_218 N_ZI_c_326_p N_SELI_c_395_n 6.45182e-19
cc_219 N_ZI_c_282_n N_SELI_c_398_n 7.64986e-19
cc_220 N_ZI_c_278_n N_SEL_c_434_n 0.00371647f
cc_221 N_ZI_c_287_n N_SEL_c_460_n 3.81736e-19
cc_222 N_ZI_XI3.X0_D N_SEL_c_438_n 9.94581e-19
cc_223 N_ZI_c_282_n N_SEL_c_438_n 0.00247421f
cc_224 N_ZI_c_280_n N_SEL_c_439_n 6.15647e-19
cc_225 N_ZI_c_326_p N_SEL_c_439_n 0.00107464f
cc_226 N_ZI_XI5.X0_D N_SEL_c_465_n 9.94581e-19
cc_227 N_ZI_c_280_n N_SEL_c_465_n 0.00243387f
cc_228 N_ZI_c_288_n N_SEL_c_453_n 0.00217047f
cc_229 N_ZI_c_282_n N_SEL_c_468_n 2.25033e-19
cc_230 N_ZI_c_278_n N_SEL_c_443_n 3.81736e-19
cc_231 N_ZI_XI6.X0_CG N_B_XI5.X0_PGS 0.00182649f
cc_232 N_Z_XI7.X0_S N_SELI_c_387_n 9.09799e-19
cc_233 Z N_SELI_c_387_n 0.00147087f
cc_234 N_SELI_c_356_n N_SEL_c_434_n 8.51271e-19
cc_235 N_SELI_c_365_n N_SEL_c_436_n 0.00269197f
cc_236 N_SELI_c_364_n N_SEL_c_438_n 0.00117605f
cc_237 N_SELI_c_356_n N_SEL_c_439_n 2.52418e-19
cc_238 N_SELI_c_364_n N_SEL_c_440_n 3.73414e-19
cc_239 N_SELI_c_365_n N_SEL_c_465_n 0.00160262f
cc_240 N_SELI_c_367_n N_SEL_c_465_n 9.78333e-19
cc_241 N_SELI_c_356_n N_SEL_c_453_n 0.00246582f
cc_242 N_SELI_c_359_n N_SEL_c_453_n 0.00269197f
cc_243 N_SELI_c_364_n N_SEL_c_468_n 2.32653e-19
cc_244 N_SELI_c_379_n N_SEL_c_468_n 3.48267e-19
cc_245 N_SELI_c_364_n N_SEL_c_442_n 9.4965e-19
cc_246 N_SELI_c_365_n N_SEL_c_442_n 2.32653e-19
cc_247 N_SELI_c_367_n N_SEL_c_442_n 3.48267e-19
cc_248 N_SELI_c_356_n N_SEL_c_443_n 9.71051e-19
cc_249 N_SELI_c_359_n N_SEL_c_443_n 6.26941e-19
cc_250 N_SELI_c_364_n N_SEL_c_444_n 3.48267e-19
cc_251 N_SELI_c_365_n N_SEL_c_444_n 7.22902e-19
cc_252 N_SELI_c_367_n N_SEL_c_444_n 0.0049864f
cc_253 N_SELI_c_379_n N_SEL_c_444_n 9.11855e-19
cc_254 N_SELI_c_364_n N_SEL_c_445_n 4.99367e-19
cc_255 N_SELI_c_365_n N_SEL_c_445_n 3.68647e-19
cc_256 N_SELI_c_367_n N_SEL_c_445_n 9.28301e-19
cc_257 N_SELI_c_379_n N_SEL_c_445_n 0.00490516f
cc_258 N_SELI_XI5.X0_CG N_B_XI5.X0_PGS 4.41254e-19
cc_259 N_SELI_c_356_n N_B_XI5.X0_PGS 2.21243e-19
cc_260 N_SELI_c_359_n N_B_XI5.X0_PGS 7.89402e-19
cc_261 N_SELI_c_367_n N_B_XI5.X0_PGS 0.00186882f
cc_262 N_SELI_c_367_n N_B_c_514_n 2.00604e-19
cc_263 N_SELI_c_371_n N_A_XI4.X0_PGS 4.65768e-19
cc_264 N_SELI_c_379_n N_A_XI4.X0_PGS 0.00276355f
cc_265 N_SELI_c_379_n N_A_c_550_n 2.00604e-19
cc_266 N_SEL_c_449_n N_B_XI5.X0_PGS 2.07014e-19
cc_267 N_SEL_c_495_p N_B_XI5.X0_PGS 4.3669e-19
cc_268 N_SEL_c_436_n N_B_XI5.X0_PGS 7.4877e-19
cc_269 N_SEL_c_443_n N_B_XI5.X0_PGS 0.00100354f
cc_270 N_SEL_c_444_n N_B_XI5.X0_PGS 0.00202689f
cc_271 N_SEL_c_468_n B 6.87706e-19
cc_272 N_SEL_c_444_n B 4.56568e-19
cc_273 N_SEL_c_495_p N_B_c_514_n 0.00234241f
cc_274 N_SEL_c_468_n N_B_c_514_n 5.02946e-19
cc_275 N_SEL_c_444_n N_B_c_514_n 0.0014909f
cc_276 N_SEL_XI4.X0_CG N_A_XI4.X0_PGS 4.54863e-19
cc_277 N_SEL_c_445_n N_A_XI4.X0_PGS 0.00276355f
cc_278 N_SEL_c_442_n A 7.05846e-19
cc_279 N_SEL_c_445_n A 4.56568e-19
cc_280 N_SEL_XI4.X0_CG N_A_c_550_n 0.00234241f
cc_281 N_SEL_c_442_n N_A_c_550_n 5.02946e-19
cc_282 N_SEL_c_445_n N_A_c_550_n 0.0014909f
cc_283 N_B_XI5.X0_PGS N_A_XI4.X0_PGS 0.00137635f
*
.ends
*
*
.subckt MUX2_HPNW4 A B S0 Y VDD VSS
xgate (VDD VSS Y S0 B A) G4_MUX2_N1_2
.ends
*
* File: G3_MUXI2_N1.pex.netlist
* Created: Wed Mar  9 13:36:32 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*







.subckt G3_MUXI2_N1_2 VSS VDD SEL B Z A
*
* A	A
* Z	Z
* B	B
* SEL	SEL
* VDD	VDD
* VSS	VSS
XI1.X0 N_SELI_XI1.X0_D N_VDD_XI1.X0_PGD N_SEL_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI2.X0 N_SELI_XI1.X0_D N_VSS_XI2.X0_PGD N_SEL_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_SELI_XI5.X0_CG N_B_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW4
XI3.X0 N_Z_XI3.X0_D N_VSS_XI3.X0_PGD N_SEL_XI3.X0_CG N_B_XI3.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI4.X0 N_Z_XI5.X0_D N_VDD_XI4.X0_PGD N_SEL_XI4.X0_CG N_A_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW4
XI0.X0 N_Z_XI3.X0_D N_VSS_XI0.X0_PGD N_SELI_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW4
*
x_PM_G3_MUXI2_N1_VSS N_VSS_XI1.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI5.X0_S N_VSS_XI3.X0_PGD N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_4_p
+ N_VSS_c_62_p N_VSS_c_21_p N_VSS_c_47_p N_VSS_c_5_p N_VSS_c_27_p N_VSS_c_18_p
+ N_VSS_c_29_p N_VSS_c_6_p N_VSS_c_20_p N_VSS_c_7_p N_VSS_c_11_p N_VSS_c_12_p
+ N_VSS_c_30_p N_VSS_c_25_p N_VSS_c_32_p N_VSS_c_37_p N_VSS_c_38_p VSS
+ N_VSS_c_13_p N_VSS_c_26_p N_VSS_c_39_p Vss PM_G3_MUXI2_N1_VSS
x_PM_G3_MUXI2_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI2.X0_S
+ N_VDD_XI5.X0_PGD N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_90_n N_VDD_c_181_p
+ N_VDD_c_91_n N_VDD_c_94_n N_VDD_c_100_n N_VDD_c_101_n N_VDD_c_107_n
+ N_VDD_c_113_n N_VDD_c_114_n N_VDD_c_117_n N_VDD_c_118_n N_VDD_c_119_n
+ N_VDD_c_120_n N_VDD_c_121_n N_VDD_c_126_n N_VDD_c_128_n VDD N_VDD_c_129_n
+ N_VDD_c_130_n N_VDD_c_135_p Vss PM_G3_MUXI2_N1_VDD
x_PM_G3_MUXI2_N1_SELI N_SELI_XI1.X0_D N_SELI_XI5.X0_CG N_SELI_XI0.X0_CG
+ N_SELI_c_188_n N_SELI_c_189_n N_SELI_c_192_n N_SELI_c_193_n N_SELI_c_209_n
+ N_SELI_c_211_n N_SELI_c_196_n N_SELI_c_198_n N_SELI_c_199_n N_SELI_c_231_p Vss
+ PM_G3_MUXI2_N1_SELI
x_PM_G3_MUXI2_N1_SEL N_SEL_XI1.X0_CG N_SEL_XI2.X0_CG N_SEL_XI3.X0_CG
+ N_SEL_XI4.X0_CG N_SEL_c_253_n N_SEL_c_254_n N_SEL_c_305_p N_SEL_c_255_n
+ N_SEL_c_257_n SEL N_SEL_c_258_n N_SEL_c_259_n N_SEL_c_274_n N_SEL_c_260_n
+ N_SEL_c_275_n N_SEL_c_262_n N_SEL_c_263_n N_SEL_c_265_n N_SEL_c_266_n Vss
+ PM_G3_MUXI2_N1_SEL
x_PM_G3_MUXI2_N1_B N_B_XI5.X0_PGS N_B_XI3.X0_PGS N_B_c_326_n N_B_c_344_n
+ N_B_c_336_n B N_B_c_328_n Vss PM_G3_MUXI2_N1_B
x_PM_G3_MUXI2_N1_Z N_Z_XI5.X0_D N_Z_XI3.X0_D N_Z_c_352_n Z Vss PM_G3_MUXI2_N1_Z
x_PM_G3_MUXI2_N1_A N_A_XI4.X0_PGS N_A_XI0.X0_PGS N_A_c_383_n A N_A_c_389_n Vss
+ PM_G3_MUXI2_N1_A
cc_1 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.0017188f
cc_2 N_VSS_XI3.X0_PGD N_VDD_XI5.X0_PGD 2.27468e-19
cc_3 N_VSS_XI0.X0_PGD N_VDD_XI4.X0_PGD 2.27468e-19
cc_4 N_VSS_c_4_p N_VDD_c_90_n 0.0017188f
cc_5 N_VSS_c_5_p N_VDD_c_91_n 9.32947e-19
cc_6 N_VSS_c_6_p N_VDD_c_91_n 3.82294e-19
cc_7 N_VSS_c_7_p N_VDD_c_91_n 4.10707e-19
cc_8 N_VSS_c_4_p N_VDD_c_94_n 2.72324e-19
cc_9 N_VSS_c_5_p N_VDD_c_94_n 0.00141228f
cc_10 N_VSS_c_6_p N_VDD_c_94_n 0.00112249f
cc_11 N_VSS_c_11_p N_VDD_c_94_n 0.00419135f
cc_12 N_VSS_c_12_p N_VDD_c_94_n 0.00124457f
cc_13 N_VSS_c_13_p N_VDD_c_94_n 7.74609e-19
cc_14 N_VSS_c_11_p N_VDD_c_100_n 0.00157719f
cc_15 N_VSS_XI2.X0_PGS N_VDD_c_101_n 2.93604e-19
cc_16 N_VSS_XI3.X0_PGD N_VDD_c_101_n 2.36238e-19
cc_17 N_VSS_c_5_p N_VDD_c_101_n 0.00181129f
cc_18 N_VSS_c_18_p N_VDD_c_101_n 7.45025e-19
cc_19 N_VSS_c_6_p N_VDD_c_101_n 9.55109e-19
cc_20 N_VSS_c_20_p N_VDD_c_101_n 2.60394e-19
cc_21 N_VSS_c_21_p N_VDD_c_107_n 0.00102426f
cc_22 N_VSS_c_18_p N_VDD_c_107_n 0.00161703f
cc_23 N_VSS_c_20_p N_VDD_c_107_n 2.03837e-19
cc_24 N_VSS_c_12_p N_VDD_c_107_n 0.0056811f
cc_25 N_VSS_c_25_p N_VDD_c_107_n 0.00454933f
cc_26 N_VSS_c_26_p N_VDD_c_107_n 7.61747e-19
cc_27 N_VSS_c_27_p N_VDD_c_113_n 0.00125492f
cc_28 N_VSS_XI4.X0_S N_VDD_c_114_n 3.7884e-19
cc_29 N_VSS_c_29_p N_VDD_c_114_n 4.73473e-19
cc_30 N_VSS_c_30_p N_VDD_c_114_n 0.00742779f
cc_31 N_VSS_c_30_p N_VDD_c_117_n 0.00149994f
cc_32 N_VSS_c_32_p N_VDD_c_118_n 4.31398e-19
cc_33 N_VSS_c_29_p N_VDD_c_119_n 2.14355e-19
cc_34 N_VSS_c_30_p N_VDD_c_120_n 0.00106317f
cc_35 N_VSS_XI4.X0_S N_VDD_c_121_n 9.5668e-19
cc_36 N_VSS_c_29_p N_VDD_c_121_n 0.00165395f
cc_37 N_VSS_c_37_p N_VDD_c_121_n 0.00364836f
cc_38 N_VSS_c_38_p N_VDD_c_121_n 0.0050309f
cc_39 N_VSS_c_39_p N_VDD_c_121_n 8.91588e-19
cc_40 N_VSS_c_18_p N_VDD_c_126_n 4.6996e-19
cc_41 N_VSS_c_38_p N_VDD_c_126_n 0.00295094f
cc_42 N_VSS_c_12_p N_VDD_c_128_n 0.00112088f
cc_43 N_VSS_c_38_p N_VDD_c_129_n 9.75645e-19
cc_44 N_VSS_c_5_p N_VDD_c_130_n 3.48267e-19
cc_45 N_VSS_c_6_p N_VDD_c_130_n 8.0279e-19
cc_46 N_VSS_XI1.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_47 N_VSS_c_47_p N_SELI_XI1.X0_D 3.48267e-19
cc_48 N_VSS_c_20_p N_SELI_c_188_n 0.00234241f
cc_49 N_VSS_XI1.X0_S N_SELI_c_189_n 3.48267e-19
cc_50 N_VSS_c_47_p N_SELI_c_189_n 8.47286e-19
cc_51 N_VSS_c_11_p N_SELI_c_189_n 2.65284e-19
cc_52 N_VSS_c_27_p N_SELI_c_192_n 0.00140233f
cc_53 N_VSS_c_18_p N_SELI_c_193_n 0.00135778f
cc_54 N_VSS_c_20_p N_SELI_c_193_n 4.99367e-19
cc_55 N_VSS_c_38_p N_SELI_c_193_n 9.07743e-19
cc_56 N_VSS_c_18_p N_SELI_c_196_n 4.56568e-19
cc_57 N_VSS_c_20_p N_SELI_c_196_n 0.0014909f
cc_58 N_VSS_c_30_p N_SELI_c_198_n 7.53578e-19
cc_59 N_VSS_c_38_p N_SELI_c_199_n 5.03655e-19
cc_60 N_VSS_XI2.X0_PGD N_SEL_c_253_n 4.12362e-19
cc_61 N_VSS_c_6_p N_SEL_c_254_n 0.00234241f
cc_62 N_VSS_c_62_p N_SEL_c_255_n 9.36847e-19
cc_63 N_VSS_c_6_p N_SEL_c_255_n 2.03369e-19
cc_64 N_VSS_c_12_p N_SEL_c_257_n 5.44326e-19
cc_65 N_VSS_c_38_p N_SEL_c_258_n 3.80099e-19
cc_66 N_VSS_c_5_p N_SEL_c_259_n 8.36018e-19
cc_67 N_VSS_c_5_p N_SEL_c_260_n 4.56568e-19
cc_68 N_VSS_c_6_p N_SEL_c_260_n 6.1245e-19
cc_69 N_VSS_c_20_p N_SEL_c_262_n 2.00604e-19
cc_70 N_VSS_c_12_p N_SEL_c_263_n 0.00127961f
cc_71 N_VSS_c_30_p N_SEL_c_263_n 2.81471e-19
cc_72 N_VSS_c_38_p N_SEL_c_265_n 4.36463e-19
cc_73 N_VSS_c_30_p N_SEL_c_266_n 0.00119312f
cc_74 N_VSS_XI2.X0_PGS N_B_c_326_n 2.96367e-19
cc_75 N_VSS_c_27_p B 0.00220388f
cc_76 N_VSS_XI5.X0_S N_B_c_328_n 0.00246958f
cc_77 N_VSS_c_27_p N_B_c_328_n 8.835e-19
cc_78 N_VSS_XI5.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_79 N_VSS_XI4.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_80 N_VSS_c_27_p N_Z_XI5.X0_D 3.48267e-19
cc_81 N_VSS_c_29_p N_Z_XI5.X0_D 3.48267e-19
cc_82 N_VSS_XI5.X0_S N_Z_c_352_n 3.48267e-19
cc_83 N_VSS_XI4.X0_S N_Z_c_352_n 3.48267e-19
cc_84 N_VSS_c_27_p N_Z_c_352_n 5.68449e-19
cc_85 N_VSS_c_29_p N_Z_c_352_n 5.69026e-19
cc_86 N_VSS_c_38_p N_Z_c_352_n 3.26224e-19
cc_87 N_VDD_XI2.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_88 N_VDD_c_94_n N_SELI_XI1.X0_D 3.7884e-19
cc_89 N_VDD_c_101_n N_SELI_XI1.X0_D 3.48267e-19
cc_90 N_VDD_c_135_p N_SELI_XI5.X0_CG 0.00237871f
cc_91 N_VDD_XI2.X0_S N_SELI_c_189_n 3.48267e-19
cc_92 N_VDD_c_94_n N_SELI_c_189_n 5.34437e-19
cc_93 N_VDD_c_101_n N_SELI_c_189_n 7.03427e-19
cc_94 N_VDD_c_94_n N_SELI_c_192_n 2.96638e-19
cc_95 N_VDD_c_121_n N_SELI_c_193_n 6.15494e-19
cc_96 N_VDD_c_113_n N_SELI_c_209_n 7.54639e-19
cc_97 N_VDD_c_135_p N_SELI_c_209_n 5.0614e-19
cc_98 N_VDD_c_113_n N_SELI_c_211_n 4.85469e-19
cc_99 N_VDD_c_135_p N_SELI_c_211_n 0.013665f
cc_100 N_VDD_c_121_n N_SELI_c_196_n 3.66936e-19
cc_101 N_VDD_c_130_n N_SEL_XI1.X0_CG 8.03148e-19
cc_102 N_VDD_XI1.X0_PGD N_SEL_c_253_n 4.25379e-19
cc_103 N_VDD_XI2.X0_S N_SEL_c_257_n 9.18655e-19
cc_104 N_VDD_c_101_n N_SEL_c_257_n 0.00161606f
cc_105 N_VDD_c_107_n N_SEL_c_258_n 2.90143e-19
cc_106 N_VDD_c_114_n N_SEL_c_258_n 3.06021e-19
cc_107 N_VDD_c_121_n N_SEL_c_258_n 6.68274e-19
cc_108 N_VDD_c_107_n N_SEL_c_274_n 2.1079e-19
cc_109 N_VDD_c_107_n N_SEL_c_275_n 2.19082e-19
cc_110 N_VDD_c_135_p N_SEL_c_275_n 2.00604e-19
cc_111 N_VDD_XI4.X0_PGD N_SEL_c_262_n 3.11814e-19
cc_112 N_VDD_c_121_n N_SEL_c_262_n 3.66936e-19
cc_113 N_VDD_c_107_n N_SEL_c_263_n 4.86613e-19
cc_114 N_VDD_c_121_n N_SEL_c_265_n 2.2501e-19
cc_115 N_VDD_c_114_n N_Z_XI5.X0_D 3.7884e-19
cc_116 N_VDD_XI2.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_117 N_VDD_XI0.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_118 N_VDD_c_101_n N_Z_XI3.X0_D 3.48267e-19
cc_119 N_VDD_c_107_n N_Z_XI3.X0_D 3.7884e-19
cc_120 N_VDD_c_119_n N_Z_XI3.X0_D 3.72199e-19
cc_121 N_VDD_XI2.X0_S N_Z_c_352_n 3.48267e-19
cc_122 N_VDD_XI0.X0_S N_Z_c_352_n 3.48267e-19
cc_123 N_VDD_c_101_n N_Z_c_352_n 8.10024e-19
cc_124 N_VDD_c_107_n N_Z_c_352_n 5.35804e-19
cc_125 N_VDD_c_114_n N_Z_c_352_n 5.35804e-19
cc_126 N_VDD_c_119_n N_Z_c_352_n 8.05266e-19
cc_127 N_VDD_c_121_n N_Z_c_352_n 7.45211e-19
cc_128 N_VDD_XI4.X0_PGD N_A_XI4.X0_PGS 0.00162178f
cc_129 N_VDD_c_121_n N_A_XI4.X0_PGS 0.0010699f
cc_130 N_VDD_c_114_n N_A_c_383_n 3.3974e-19
cc_131 N_VDD_c_121_n N_A_c_383_n 4.15738e-19
cc_132 N_VDD_c_113_n A 5.43314e-19
cc_133 N_VDD_c_114_n A 0.00141439f
cc_134 N_VDD_c_121_n A 5.04211e-19
cc_135 N_VDD_c_135_p A 3.48267e-19
cc_136 N_VDD_c_181_p N_A_c_389_n 0.00480616f
cc_137 N_VDD_c_113_n N_A_c_389_n 3.89161e-19
cc_138 N_VDD_c_114_n N_A_c_389_n 0.00117371f
cc_139 N_VDD_c_121_n N_A_c_389_n 4.41003e-19
cc_140 N_VDD_c_135_p N_A_c_389_n 6.39485e-19
cc_141 N_SELI_c_189_n N_SEL_c_253_n 8.93041e-19
cc_142 N_SELI_c_192_n N_SEL_c_253_n 3.46631e-19
cc_143 N_SELI_c_209_n N_SEL_c_257_n 0.00339809f
cc_144 N_SELI_c_193_n N_SEL_c_258_n 0.00240446f
cc_145 N_SELI_c_189_n N_SEL_c_259_n 0.0021504f
cc_146 N_SELI_c_192_n N_SEL_c_259_n 0.00339809f
cc_147 N_SELI_c_189_n N_SEL_c_260_n 9.71051e-19
cc_148 N_SELI_c_192_n N_SEL_c_260_n 6.41327e-19
cc_149 N_SELI_c_209_n N_SEL_c_275_n 7.09664e-19
cc_150 N_SELI_c_211_n N_SEL_c_275_n 0.00496695f
cc_151 N_SELI_c_196_n N_SEL_c_275_n 8.74049e-19
cc_152 N_SELI_c_193_n N_SEL_c_262_n 4.99367e-19
cc_153 N_SELI_c_211_n N_SEL_c_262_n 8.86313e-19
cc_154 N_SELI_c_196_n N_SEL_c_262_n 0.00491002f
cc_155 N_SELI_c_193_n N_SEL_c_263_n 0.00165721f
cc_156 N_SELI_c_209_n N_SEL_c_263_n 4.70859e-19
cc_157 N_SELI_c_198_n N_SEL_c_263_n 9.36901e-19
cc_158 N_SELI_c_231_p N_SEL_c_263_n 7.85443e-19
cc_159 N_SELI_c_189_n N_SEL_c_265_n 2.46723e-19
cc_160 N_SELI_c_209_n N_SEL_c_265_n 2.46502e-19
cc_161 N_SELI_c_199_n N_SEL_c_265_n 0.00142585f
cc_162 N_SELI_c_209_n N_SEL_c_266_n 0.00166116f
cc_163 N_SELI_c_198_n N_SEL_c_266_n 7.57935e-19
cc_164 N_SELI_XI5.X0_CG N_B_XI5.X0_PGS 4.34645e-19
cc_165 N_SELI_c_211_n N_B_XI5.X0_PGS 6.90642e-19
cc_166 N_SELI_c_189_n N_B_XI3.X0_PGS 2.37944e-19
cc_167 N_SELI_c_192_n N_B_XI3.X0_PGS 3.60699e-19
cc_168 N_SELI_c_211_n N_B_XI3.X0_PGS 5.45575e-19
cc_169 N_SELI_c_192_n N_B_c_326_n 3.87281e-19
cc_170 N_SELI_c_192_n N_B_c_336_n 5.40503e-19
cc_171 N_SELI_c_192_n B 0.0012892f
cc_172 N_SELI_c_192_n N_B_c_328_n 0.00106294f
cc_173 N_SELI_c_189_n N_Z_c_352_n 5.41397e-19
cc_174 N_SELI_c_193_n N_Z_c_352_n 0.00205681f
cc_175 N_SELI_c_209_n N_Z_c_352_n 0.00246976f
cc_176 N_SELI_c_211_n N_Z_c_352_n 9.16045e-19
cc_177 N_SELI_c_188_n N_A_XI4.X0_PGS 4.5346e-19
cc_178 N_SELI_c_196_n N_A_XI4.X0_PGS 0.00276355f
cc_179 N_SELI_c_196_n N_A_c_389_n 2.00604e-19
cc_180 N_SEL_c_254_n N_B_XI3.X0_PGS 2.04953e-19
cc_181 N_SEL_c_305_p N_B_XI3.X0_PGS 4.64062e-19
cc_182 N_SEL_c_257_n N_B_XI3.X0_PGS 8.04174e-19
cc_183 N_SEL_c_260_n N_B_XI3.X0_PGS 0.00100354f
cc_184 N_SEL_c_275_n N_B_XI3.X0_PGS 0.00142122f
cc_185 N_SEL_c_257_n N_B_c_344_n 2.97958e-19
cc_186 N_SEL_c_260_n N_B_c_344_n 3.50453e-19
cc_187 N_SEL_c_260_n N_B_c_328_n 9.99041e-19
cc_188 N_SEL_c_258_n N_Z_c_352_n 0.00187327f
cc_189 N_SEL_c_274_n N_Z_c_352_n 0.00194252f
cc_190 N_SEL_c_275_n N_Z_c_352_n 9.12105e-19
cc_191 N_SEL_c_262_n N_Z_c_352_n 9.02042e-19
cc_192 N_SEL_c_263_n N_Z_c_352_n 8.60225e-19
cc_193 N_SEL_c_265_n N_Z_c_352_n 0.0021646f
cc_194 N_SEL_c_266_n N_Z_c_352_n 8.38981e-19
cc_195 N_SEL_XI4.X0_CG N_A_XI4.X0_PGS 4.42555e-19
cc_196 N_SEL_c_262_n N_A_XI4.X0_PGS 0.00276355f
cc_197 N_SEL_c_258_n A 7.0885e-19
cc_198 N_SEL_c_262_n A 4.56568e-19
cc_199 N_SEL_XI4.X0_CG N_A_c_389_n 0.00234241f
cc_200 N_SEL_c_258_n N_A_c_389_n 4.99367e-19
cc_201 N_SEL_c_262_n N_A_c_389_n 0.0014909f
cc_202 N_B_XI5.X0_PGS N_A_XI4.X0_PGS 0.00137535f
*
.ends
*
*
.subckt MUXI2_HPNW4 A B S0 Y VDD VSS
xgate (VSS VDD S0 B Y A) G3_MUXI2_N1_2
.ends
*
* File: G2_NAND2_N1.pex.netlist
* Created: Tue Feb 22 16:31:07 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*





.subckt G2_NAND2_N1_2 VSS VDD A Z B
*
* B	B
* Z	Z
* A	A
* VDD	VDD
* VSS	VSS
XI7.X0 N_Z_XI7.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_B_XI7.X0_PGS N_VSS_XI7.X0_S
+ TIGFET_HPNW4
XI8.X0 N_Z_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI9.X0 N_Z_XI8.X0_D N_VSS_XI9.X0_PGD N_B_XI9.X0_CG N_VSS_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW4
*
x_PM_G2_NAND2_N1_VSS N_VSS_XI7.X0_S N_VSS_XI8.X0_PGD N_VSS_XI8.X0_PGS
+ N_VSS_XI9.X0_PGD N_VSS_XI9.X0_PGS N_VSS_c_6_p N_VSS_c_18_p N_VSS_c_1_p
+ N_VSS_c_4_p N_VSS_c_5_p VSS N_VSS_c_9_p N_VSS_c_10_p Vss PM_G2_NAND2_N1_VSS
x_PM_G2_NAND2_N1_VDD N_VDD_XI7.X0_PGD N_VDD_XI8.X0_S N_VDD_XI9.X0_S N_VDD_c_61_p
+ N_VDD_c_54_p N_VDD_c_29_n N_VDD_c_33_n N_VDD_c_37_n N_VDD_c_57_p N_VDD_c_38_n
+ VDD N_VDD_c_43_p Vss PM_G2_NAND2_N1_VDD
x_PM_G2_NAND2_N1_A N_A_XI7.X0_CG N_A_XI8.X0_CG N_A_c_71_n N_A_c_72_n A
+ N_A_c_79_n N_A_c_75_n Vss PM_G2_NAND2_N1_A
x_PM_G2_NAND2_N1_Z N_Z_XI7.X0_D N_Z_XI8.X0_D N_Z_c_94_n Z Vss PM_G2_NAND2_N1_Z
x_PM_G2_NAND2_N1_B N_B_XI7.X0_PGS N_B_XI9.X0_CG N_B_c_117_n N_B_c_119_n
+ N_B_c_123_n N_B_c_127_n B Vss PM_G2_NAND2_N1_B
cc_1 N_VSS_c_1_p N_VDD_XI8.X0_S 0.00136022f
cc_2 N_VSS_XI8.X0_PGS N_VDD_c_29_n 4.05134e-19
cc_3 N_VSS_c_1_p N_VDD_c_29_n 0.00385472f
cc_4 N_VSS_c_4_p N_VDD_c_29_n 0.00232594f
cc_5 N_VSS_c_5_p N_VDD_c_29_n 0.00101015f
cc_6 N_VSS_c_6_p N_VDD_c_33_n 0.00171596f
cc_7 N_VSS_c_4_p N_VDD_c_33_n 0.00161703f
cc_8 N_VSS_c_5_p N_VDD_c_33_n 2.03837e-19
cc_9 N_VSS_c_9_p N_VDD_c_33_n 0.00286543f
cc_10 N_VSS_c_10_p N_VDD_c_37_n 0.00103397f
cc_11 N_VSS_XI9.X0_PGS N_VDD_c_38_n 4.47716e-19
cc_12 N_VSS_c_1_p N_VDD_c_38_n 2.23518e-19
cc_13 N_VSS_c_4_p N_VDD_c_38_n 5.24284e-19
cc_14 N_VSS_c_5_p N_A_c_71_n 0.00234241f
cc_15 N_VSS_c_1_p N_A_c_72_n 0.00297841f
cc_16 N_VSS_c_4_p N_A_c_72_n 8.12473e-19
cc_17 N_VSS_c_5_p N_A_c_72_n 5.42695e-19
cc_18 N_VSS_c_18_p N_A_c_75_n 7.84334e-19
cc_19 N_VSS_c_4_p N_A_c_75_n 4.56568e-19
cc_20 N_VSS_c_5_p N_A_c_75_n 0.00184767f
cc_21 N_VSS_XI7.X0_S N_Z_XI7.X0_D 3.43419e-19
cc_22 N_VSS_c_1_p N_Z_XI7.X0_D 3.48267e-19
cc_23 N_VSS_XI7.X0_S N_Z_c_94_n 3.48267e-19
cc_24 N_VSS_c_1_p N_Z_c_94_n 0.00178967f
cc_25 N_VSS_XI8.X0_PGD N_B_c_117_n 6.72196e-19
cc_26 N_VSS_XI9.X0_PGD N_B_c_117_n 6.72196e-19
cc_27 N_VSS_XI8.X0_PGS N_B_c_119_n 7.91098e-19
cc_28 N_VDD_XI7.X0_PGD N_A_XI7.X0_CG 4.91184e-19
cc_29 N_VDD_XI7.X0_PGD N_A_c_79_n 2.88617e-19
cc_30 N_VDD_c_43_p N_A_c_79_n 7.96439e-19
cc_31 N_VDD_c_33_n N_A_c_75_n 2.29043e-19
cc_32 N_VDD_c_43_p N_Z_XI7.X0_D 0.00132057f
cc_33 N_VDD_XI8.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_34 N_VDD_XI9.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_35 N_VDD_c_29_n N_Z_XI8.X0_D 3.48267e-19
cc_36 N_VDD_c_33_n N_Z_XI8.X0_D 3.7884e-19
cc_37 N_VDD_c_38_n N_Z_XI8.X0_D 3.48267e-19
cc_38 N_VDD_XI7.X0_PGD N_Z_c_94_n 3.00781e-19
cc_39 N_VDD_XI8.X0_S N_Z_c_94_n 3.48267e-19
cc_40 N_VDD_XI9.X0_S N_Z_c_94_n 3.48267e-19
cc_41 N_VDD_c_54_p N_Z_c_94_n 7.07078e-19
cc_42 N_VDD_c_29_n N_Z_c_94_n 5.69026e-19
cc_43 N_VDD_c_33_n N_Z_c_94_n 7.07375e-19
cc_44 N_VDD_c_57_p N_Z_c_94_n 0.00174191f
cc_45 N_VDD_c_38_n N_Z_c_94_n 0.00291831f
cc_46 N_VDD_c_43_p N_Z_c_94_n 8.835e-19
cc_47 N_VDD_XI7.X0_PGD N_B_XI7.X0_PGS 0.00320747f
cc_48 N_VDD_c_61_p N_B_c_117_n 0.0097987f
cc_49 N_VDD_c_38_n N_B_c_117_n 2.48119e-19
cc_50 N_VDD_c_33_n N_B_c_123_n 4.73957e-19
cc_51 N_VDD_c_57_p N_B_c_123_n 3.81676e-19
cc_52 N_VDD_c_38_n N_B_c_123_n 0.001001f
cc_53 N_VDD_c_43_p N_B_c_123_n 0.00150149f
cc_54 N_VDD_c_33_n N_B_c_127_n 4.10393e-19
cc_55 N_VDD_c_57_p N_B_c_127_n 5.19718e-19
cc_56 N_VDD_c_38_n N_B_c_127_n 0.00144738f
cc_57 N_VDD_c_43_p N_B_c_127_n 3.81676e-19
cc_58 N_A_c_72_n N_Z_c_94_n 0.00754545f
cc_59 N_A_c_79_n N_Z_c_94_n 9.58524e-19
cc_60 N_A_c_75_n N_Z_c_94_n 9.18163e-19
cc_61 N_A_XI7.X0_CG N_B_XI7.X0_PGS 4.5346e-19
cc_62 N_A_c_72_n N_B_XI7.X0_PGS 2.82086e-19
cc_63 N_A_c_79_n N_B_XI7.X0_PGS 5.70584e-19
cc_64 N_A_c_72_n N_B_c_117_n 3.21972e-19
cc_65 N_A_c_79_n N_B_c_117_n 0.0014179f
cc_66 N_A_c_75_n N_B_c_117_n 0.00112482f
cc_67 N_A_c_75_n N_B_c_123_n 9.27569e-19
cc_68 N_Z_c_94_n N_B_c_117_n 3.90525e-19
cc_69 N_Z_c_94_n N_B_c_123_n 9.49424e-19
cc_70 N_Z_c_94_n N_B_c_127_n 0.00147334f
*
.ends
*
*
.subckt NAND2_HPNW4 A B Y VDD VSS
xgate (VSS VDD A Y B) G2_NAND2_N1_2
.ends
*
* File: G2_NOR2_N1.pex.netlist
* Created: Mon Feb 28 09:28:35 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*





.subckt G2_NOR2_N1_2 VSS VDD B Z A
*
* A	A
* Z	Z
* B	B
* VDD	VDD
* VSS	VSS
XI2.X0 N_Z_XI2.X0_D N_VDD_XI2.X0_PGD N_B_XI2.X0_CG N_VDD_XI2.X0_PGS
+ N_VSS_XI2.X0_S TIGFET_HPNW4
XI0.X0 N_Z_XI0.X0_D N_VSS_XI0.X0_PGD N_B_XI0.X0_CG N_A_XI0.X0_PGS N_VDD_XI0.X0_S
+ TIGFET_HPNW4
XI1.X0 N_Z_XI0.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
*
x_PM_G2_NOR2_N1_VSS N_VSS_XI2.X0_S N_VSS_XI0.X0_PGD N_VSS_XI1.X0_S N_VSS_c_31_p
+ N_VSS_c_2_p N_VSS_c_4_p N_VSS_c_7_p N_VSS_c_37_p N_VSS_c_8_p VSS N_VSS_c_6_p
+ N_VSS_c_16_p N_VSS_c_19_p N_VSS_c_17_p N_VSS_c_22_p N_VSS_c_18_p Vss
+ PM_G2_NOR2_N1_VSS
x_PM_G2_NOR2_N1_VDD N_VDD_XI2.X0_PGD N_VDD_XI2.X0_PGS N_VDD_XI0.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_c_45_n N_VDD_c_90_p N_VDD_c_46_n
+ N_VDD_c_50_n N_VDD_c_53_n N_VDD_c_55_n N_VDD_c_56_n N_VDD_c_62_n VDD
+ N_VDD_c_72_p N_VDD_c_63_n N_VDD_c_66_n N_VDD_c_69_p N_VDD_c_67_n Vss
+ PM_G2_NOR2_N1_VDD
x_PM_G2_NOR2_N1_B N_B_XI2.X0_CG N_B_XI0.X0_CG N_B_c_104_n N_B_c_95_n N_B_c_96_n
+ B N_B_c_99_n N_B_c_100_n Vss PM_G2_NOR2_N1_B
x_PM_G2_NOR2_N1_Z N_Z_XI2.X0_D N_Z_XI0.X0_D N_Z_c_124_n Z Vss PM_G2_NOR2_N1_Z
x_PM_G2_NOR2_N1_A N_A_XI0.X0_PGS N_A_XI1.X0_CG N_A_c_141_n N_A_c_145_n
+ N_A_c_147_n A Vss PM_G2_NOR2_N1_A
cc_1 N_VSS_XI0.X0_PGD N_VDD_XI1.X0_PGD 0.00180308f
cc_2 N_VSS_c_2_p N_VDD_c_45_n 0.00180308f
cc_3 N_VSS_XI2.X0_S N_VDD_c_46_n 9.5668e-19
cc_4 N_VSS_c_4_p N_VDD_c_46_n 0.00165395f
cc_5 VSS N_VDD_c_46_n 0.00476397f
cc_6 N_VSS_c_6_p N_VDD_c_46_n 0.00186257f
cc_7 N_VSS_c_7_p N_VDD_c_50_n 4.43871e-19
cc_8 N_VSS_c_8_p N_VDD_c_50_n 3.66936e-19
cc_9 VSS N_VDD_c_50_n 0.00285866f
cc_10 N_VSS_XI2.X0_S N_VDD_c_53_n 3.7884e-19
cc_11 N_VSS_c_4_p N_VDD_c_53_n 0.00104703f
cc_12 N_VSS_c_4_p N_VDD_c_55_n 7.47067e-19
cc_13 N_VSS_c_2_p N_VDD_c_56_n 3.37151e-19
cc_14 N_VSS_c_7_p N_VDD_c_56_n 0.00141228f
cc_15 N_VSS_c_8_p N_VDD_c_56_n 0.00112249f
cc_16 N_VSS_c_16_p N_VDD_c_56_n 0.0034844f
cc_17 N_VSS_c_17_p N_VDD_c_56_n 0.00588723f
cc_18 N_VSS_c_18_p N_VDD_c_56_n 7.74609e-19
cc_19 N_VSS_c_19_p N_VDD_c_62_n 0.00106075f
cc_20 N_VSS_c_7_p N_VDD_c_63_n 0.00106112f
cc_21 N_VSS_c_8_p N_VDD_c_63_n 3.95933e-19
cc_22 N_VSS_c_22_p N_VDD_c_63_n 3.86251e-19
cc_23 VSS N_VDD_c_66_n 0.00116512f
cc_24 N_VSS_c_7_p N_VDD_c_67_n 3.44698e-19
cc_25 N_VSS_c_8_p N_VDD_c_67_n 7.95135e-19
cc_26 N_VSS_c_8_p N_B_c_95_n 0.00234321f
cc_27 N_VSS_c_7_p N_B_c_96_n 8.39582e-19
cc_28 N_VSS_c_8_p N_B_c_96_n 5.42695e-19
cc_29 VSS N_B_c_96_n 0.00148607f
cc_30 N_VSS_c_8_p N_B_c_99_n 2.00604e-19
cc_31 N_VSS_c_31_p N_B_c_100_n 8.37306e-19
cc_32 N_VSS_c_7_p N_B_c_100_n 4.56568e-19
cc_33 N_VSS_c_8_p N_B_c_100_n 0.00173573f
cc_34 N_VSS_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_35 N_VSS_c_4_p N_Z_XI2.X0_D 3.48267e-19
cc_36 N_VSS_XI1.X0_S N_Z_XI0.X0_D 3.43419e-19
cc_37 N_VSS_c_37_p N_Z_XI0.X0_D 3.48267e-19
cc_38 N_VSS_c_4_p N_Z_c_124_n 8.89782e-19
cc_39 N_VSS_c_37_p N_Z_c_124_n 6.0686e-19
cc_40 VSS N_Z_c_124_n 4.63431e-19
cc_41 N_VSS_c_17_p N_Z_c_124_n 2.55365e-19
cc_42 N_VSS_XI0.X0_PGD N_A_c_141_n 9.39677e-19
cc_43 N_VSS_c_2_p N_A_c_141_n 2.16729e-19
cc_44 N_VDD_c_69_p N_B_XI2.X0_CG 0.00237871f
cc_45 N_VDD_c_69_p N_B_c_104_n 0.0010681f
cc_46 N_VDD_c_46_n N_B_c_96_n 0.0025037f
cc_47 N_VDD_c_72_p N_B_c_96_n 7.41679e-19
cc_48 N_VDD_c_69_p N_B_c_96_n 5.48133e-19
cc_49 N_VDD_c_46_n N_B_c_99_n 4.9897e-19
cc_50 N_VDD_c_72_p N_B_c_99_n 4.91501e-19
cc_51 N_VDD_c_69_p N_B_c_99_n 0.00150793f
cc_52 N_VDD_c_46_n N_B_c_100_n 3.66936e-19
cc_53 N_VDD_c_69_p N_B_c_100_n 2.00604e-19
cc_54 N_VDD_XI0.X0_S N_Z_XI0.X0_D 3.43419e-19
cc_55 N_VDD_c_55_n N_Z_XI0.X0_D 3.72199e-19
cc_56 N_VDD_c_56_n N_Z_XI0.X0_D 3.7884e-19
cc_57 N_VDD_XI0.X0_S N_Z_c_124_n 3.48267e-19
cc_58 N_VDD_c_46_n N_Z_c_124_n 5.1034e-19
cc_59 N_VDD_c_55_n N_Z_c_124_n 7.89245e-19
cc_60 N_VDD_c_56_n N_Z_c_124_n 5.36364e-19
cc_61 N_VDD_XI2.X0_PGD N_A_c_141_n 5.10213e-19
cc_62 N_VDD_XI1.X0_PGD N_A_c_141_n 2.48727e-19
cc_63 N_VDD_XI2.X0_PGS N_A_c_145_n 6.4837e-19
cc_64 N_VDD_c_46_n N_A_c_145_n 3.16598e-19
cc_65 N_VDD_c_90_p N_A_c_147_n 8.9931e-19
cc_66 N_VDD_c_63_n N_A_c_147_n 4.91217e-19
cc_67 N_VDD_c_67_n N_A_c_147_n 0.00320668f
cc_68 N_VDD_c_63_n A 6.1931e-19
cc_69 N_VDD_c_67_n A 4.56568e-19
cc_70 N_B_c_96_n N_Z_c_124_n 0.00744925f
cc_71 N_B_c_99_n N_Z_c_124_n 9.58524e-19
cc_72 N_B_c_100_n N_Z_c_124_n 8.92526e-19
cc_73 N_B_c_95_n N_A_XI0.X0_PGS 4.5346e-19
cc_74 N_B_c_100_n N_A_XI0.X0_PGS 7.86826e-19
cc_75 N_B_c_99_n N_A_c_141_n 9.25308e-19
cc_76 N_B_c_100_n N_A_c_147_n 7.50183e-19
cc_77 N_Z_c_124_n N_A_c_141_n 9.72643e-19
cc_78 N_Z_c_124_n N_A_c_147_n 9.67259e-19
cc_79 N_Z_c_124_n A 0.00155484f
*
.ends
*
*
.subckt NOR2_HPNW4 A B Y VDD VSS
xgate (VSS VDD B Y A) G2_NOR2_N1_2
.ends
*
* File: G2_OAI21_N1.pex.netlist
* Created: Wed Feb 23 15:42:41 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*






.subckt G2_OAI21_N1_2 VSS VDD B A Z C
*
* C	C
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI1.X0 N_Z_XI1.X0_D N_VDD_XI1.X0_PGD N_B_XI1.X0_CG N_C_XI1.X0_PGS N_VSS_XI1.X0_S
+ TIGFET_HPNW4
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_A_XI6.X0_PGS N_VDD_XI6.X0_S
+ TIGFET_HPNW4
XI5.X0 N_Z_XI1.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_C_XI5.X0_PGS N_VSS_XI5.X0_S
+ TIGFET_HPNW4
XI7.X0 N_Z_XI6.X0_D N_VSS_XI7.X0_PGD N_C_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW4
*
x_PM_G2_OAI21_N1_VSS N_VSS_XI1.X0_S N_VSS_XI6.X0_PGD N_VSS_XI5.X0_S
+ N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS N_VSS_c_22_p N_VSS_c_44_p N_VSS_c_1_p
+ N_VSS_c_23_p N_VSS_c_9_p N_VSS_c_24_p N_VSS_c_2_p N_VSS_c_3_p N_VSS_c_7_p
+ N_VSS_c_12_p N_VSS_c_10_p N_VSS_c_16_p VSS Vss PM_G2_OAI21_N1_VSS
x_PM_G2_OAI21_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI6.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI7.X0_S N_VDD_c_50_n N_VDD_c_53_n N_VDD_c_54_n N_VDD_c_55_n
+ N_VDD_c_75_p N_VDD_c_57_n N_VDD_c_60_n N_VDD_c_63_n VDD N_VDD_c_72_p Vss
+ PM_G2_OAI21_N1_VDD
x_PM_G2_OAI21_N1_B N_B_XI1.X0_CG N_B_XI6.X0_CG N_B_c_102_n N_B_c_109_p
+ N_B_c_101_n B N_B_c_105_n N_B_c_107_n Vss PM_G2_OAI21_N1_B
x_PM_G2_OAI21_N1_A N_A_XI6.X0_PGS N_A_XI5.X0_CG N_A_c_139_n N_A_c_149_n
+ N_A_c_125_n N_A_c_127_n N_A_c_131_n A N_A_c_137_n Vss PM_G2_OAI21_N1_A
x_PM_G2_OAI21_N1_Z N_Z_XI1.X0_D N_Z_XI6.X0_D N_Z_c_171_n Z Vss PM_G2_OAI21_N1_Z
x_PM_G2_OAI21_N1_C N_C_XI1.X0_PGS N_C_XI5.X0_PGS N_C_XI7.X0_CG N_C_c_197_n
+ N_C_c_219_n N_C_c_199_n N_C_c_202_n N_C_c_203_n C Vss PM_G2_OAI21_N1_C
cc_1 N_VSS_c_1_p N_VDD_c_50_n 0.00187494f
cc_2 N_VSS_c_2_p N_VDD_c_50_n 0.00510452f
cc_3 N_VSS_c_3_p N_VDD_c_50_n 0.00186257f
cc_4 N_VSS_c_1_p N_VDD_c_53_n 0.0010904f
cc_5 N_VSS_c_2_p N_VDD_c_54_n 0.0014876f
cc_6 N_VSS_c_1_p N_VDD_c_55_n 7.48363e-19
cc_7 N_VSS_c_7_p N_VDD_c_55_n 4.59722e-19
cc_8 N_VSS_XI5.X0_S N_VDD_c_57_n 3.7884e-19
cc_9 N_VSS_c_9_p N_VDD_c_57_n 5.11058e-19
cc_10 N_VSS_c_10_p N_VDD_c_57_n 5.35974e-19
cc_11 N_VSS_c_9_p N_VDD_c_60_n 2.14355e-19
cc_12 N_VSS_c_12_p N_VDD_c_60_n 4.59722e-19
cc_13 N_VSS_c_10_p N_VDD_c_60_n 5.34009e-19
cc_14 N_VSS_c_9_p N_VDD_c_63_n 0.00187494f
cc_15 N_VSS_c_10_p N_VDD_c_63_n 0.00186257f
cc_16 N_VSS_c_16_p N_VDD_c_63_n 0.00730042f
cc_17 N_VSS_c_2_p N_B_c_101_n 5.86846e-19
cc_18 N_VSS_XI6.X0_PGD N_A_XI6.X0_PGS 0.00164631f
cc_19 N_VSS_c_7_p N_A_c_125_n 8.83597e-19
cc_20 N_VSS_c_16_p N_A_c_125_n 4.02032e-19
cc_21 N_VSS_XI6.X0_PGD N_A_c_127_n 3.11814e-19
cc_22 N_VSS_c_22_p N_A_c_127_n 0.00322564f
cc_23 N_VSS_c_23_p N_A_c_127_n 3.44698e-19
cc_24 N_VSS_c_24_p N_A_c_127_n 6.61253e-19
cc_25 N_VSS_c_24_p N_A_c_131_n 3.77503e-19
cc_26 N_VSS_c_23_p A 8.59446e-19
cc_27 N_VSS_c_24_p A 3.44698e-19
cc_28 N_VSS_c_2_p A 0.00272781f
cc_29 N_VSS_c_7_p A 0.00211023f
cc_30 N_VSS_c_16_p A 0.00133784f
cc_31 N_VSS_c_2_p N_A_c_137_n 0.00291082f
cc_32 N_VSS_XI1.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_33 N_VSS_XI5.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_34 N_VSS_c_1_p N_Z_XI1.X0_D 3.48267e-19
cc_35 N_VSS_c_9_p N_Z_XI1.X0_D 3.48267e-19
cc_36 N_VSS_XI1.X0_S N_Z_c_171_n 3.48267e-19
cc_37 N_VSS_XI5.X0_S N_Z_c_171_n 3.48267e-19
cc_38 N_VSS_c_1_p N_Z_c_171_n 5.69026e-19
cc_39 N_VSS_c_9_p N_Z_c_171_n 5.69026e-19
cc_40 N_VSS_c_7_p N_Z_c_171_n 4.84633e-19
cc_41 N_VSS_c_16_p N_Z_c_171_n 4.50981e-19
cc_42 N_VSS_XI6.X0_PGD N_C_c_197_n 6.77138e-19
cc_43 N_VSS_XI7.X0_PGD N_C_c_197_n 6.77138e-19
cc_44 N_VSS_c_44_p N_C_c_199_n 8.9608e-19
cc_45 N_VSS_c_23_p N_C_c_199_n 4.56568e-19
cc_46 N_VSS_c_24_p N_C_c_199_n 0.00315719f
cc_47 N_VSS_XI7.X0_PGS N_C_c_202_n 7.91098e-19
cc_48 N_VSS_c_23_p N_C_c_203_n 5.37794e-19
cc_49 N_VSS_c_24_p N_C_c_203_n 4.56568e-19
cc_50 N_VDD_c_53_n N_B_c_102_n 2.44914e-19
cc_51 N_VDD_c_50_n N_B_c_101_n 0.00216638f
cc_52 N_VDD_c_53_n N_B_c_101_n 2.85486e-19
cc_53 N_VDD_c_50_n N_B_c_105_n 3.66936e-19
cc_54 N_VDD_c_53_n N_B_c_105_n 2.29043e-19
cc_55 N_VDD_c_50_n N_B_c_107_n 4.1997e-19
cc_56 N_VDD_c_72_p N_A_XI5.X0_CG 0.00237871f
cc_57 N_VDD_c_72_p N_A_c_139_n 0.00106215f
cc_58 N_VDD_c_53_n N_A_c_125_n 9.72202e-19
cc_59 N_VDD_c_75_p N_A_c_125_n 7.80108e-19
cc_60 N_VDD_c_63_n N_A_c_125_n 6.23587e-19
cc_61 N_VDD_c_72_p N_A_c_125_n 4.87728e-19
cc_62 N_VDD_c_75_p N_A_c_131_n 4.85469e-19
cc_63 N_VDD_c_63_n N_A_c_131_n 3.66936e-19
cc_64 N_VDD_c_72_p N_A_c_131_n 0.0014909f
cc_65 N_VDD_c_50_n N_A_c_137_n 6.23756e-19
cc_66 N_VDD_c_53_n N_A_c_137_n 2.0345e-19
cc_67 N_VDD_c_53_n N_Z_XI1.X0_D 3.7884e-19
cc_68 N_VDD_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_69 N_VDD_XI7.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_70 N_VDD_c_55_n N_Z_XI6.X0_D 3.72199e-19
cc_71 N_VDD_c_60_n N_Z_XI6.X0_D 3.72199e-19
cc_72 N_VDD_XI6.X0_S N_Z_c_171_n 3.48267e-19
cc_73 N_VDD_XI7.X0_S N_Z_c_171_n 3.48267e-19
cc_74 N_VDD_c_50_n N_Z_c_171_n 3.87755e-19
cc_75 N_VDD_c_53_n N_Z_c_171_n 6.81554e-19
cc_76 N_VDD_c_55_n N_Z_c_171_n 5.6271e-19
cc_77 N_VDD_c_60_n N_Z_c_171_n 7.76033e-19
cc_78 N_VDD_c_63_n N_Z_c_171_n 0.0010014f
cc_79 N_VDD_c_50_n N_C_XI1.X0_PGS 6.09123e-19
cc_80 N_VDD_c_63_n N_C_XI5.X0_PGS 6.28572e-19
cc_81 N_VDD_XI1.X0_PGD N_C_c_197_n 6.72196e-19
cc_82 N_VDD_XI5.X0_PGD N_C_c_197_n 6.76891e-19
cc_83 N_VDD_c_63_n N_C_c_199_n 4.79801e-19
cc_84 N_VDD_c_63_n N_C_c_203_n 3.46645e-19
cc_85 N_B_c_107_n N_A_c_149_n 8.43061e-19
cc_86 N_B_c_109_p N_A_c_127_n 0.00234241f
cc_87 N_B_c_101_n N_A_c_127_n 5.28799e-19
cc_88 N_B_c_107_n N_A_c_127_n 0.00173494f
cc_89 N_B_c_105_n N_A_c_131_n 8.86454e-19
cc_90 N_B_c_101_n A 0.00306515f
cc_91 N_B_c_107_n A 4.56568e-19
cc_92 N_B_c_101_n N_A_c_137_n 6.59436e-19
cc_93 N_B_c_101_n N_Z_c_171_n 0.00673203f
cc_94 N_B_c_105_n N_Z_c_171_n 9.17696e-19
cc_95 N_B_c_107_n N_Z_c_171_n 9.18163e-19
cc_96 N_B_XI1.X0_CG N_C_XI1.X0_PGS 4.42555e-19
cc_97 N_B_c_105_n N_C_XI1.X0_PGS 0.001089f
cc_98 N_B_c_105_n N_C_c_197_n 6.02551e-19
cc_99 N_B_c_107_n N_C_c_197_n 0.00107456f
cc_100 N_B_c_107_n N_C_c_199_n 9.3196e-19
cc_101 N_A_c_125_n N_Z_c_171_n 0.00382179f
cc_102 A N_Z_c_171_n 0.00134325f
cc_103 N_A_XI5.X0_CG N_C_XI5.X0_PGS 4.42555e-19
cc_104 N_A_c_131_n N_C_XI5.X0_PGS 0.001089f
cc_105 N_A_c_131_n N_C_c_197_n 6.59241e-19
cc_106 N_A_XI6.X0_PGS N_C_c_219_n 7.91098e-19
cc_107 N_A_c_125_n N_C_c_199_n 5.38228e-19
cc_108 N_A_c_127_n N_C_c_199_n 2.62413e-19
cc_109 N_A_c_131_n N_C_c_199_n 0.0021499f
cc_110 N_A_c_125_n N_C_c_203_n 8.10255e-19
cc_111 N_Z_c_171_n N_C_c_197_n 4.9701e-19
cc_112 N_Z_c_171_n N_C_c_199_n 9.61365e-19
cc_113 N_Z_c_171_n N_C_c_203_n 0.00143964f
*
.ends
*
*
.subckt OAI21_HPNW4 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 A0 Y B0) G2_OAI21_N1_2
.ends
*
* File: G3_OR2_N1.pex.netlist
* Created: Tue Mar  1 11:26:38 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*






.subckt G3_OR2_N1_2 VSS VDD B A Z
*
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI2.X0 N_NET21_XI2.X0_D N_VDD_XI2.X0_PGD N_B_XI2.X0_CG N_VDD_XI2.X0_PGS
+ N_VSS_XI2.X0_S TIGFET_HPNW4
XI0.X0 N_NET21_XI0.X0_D N_VSS_XI0.X0_PGD N_B_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW4
XI1.X0 N_NET21_XI0.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_NET21_XI3.X0_CG N_VDD_XI3.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI4.X0 N_Z_XI3.X0_D N_VSS_XI4.X0_PGD N_NET21_XI4.X0_CG N_VSS_XI4.X0_PGS
+ N_VDD_XI4.X0_S TIGFET_HPNW4
*
x_PM_G3_OR2_N1_VSS N_VSS_XI2.X0_S N_VSS_XI0.X0_PGD N_VSS_XI1.X0_S
+ N_VSS_XI4.X0_PGD N_VSS_XI4.X0_PGS N_VSS_c_32_p N_VSS_c_4_p N_VSS_c_51_p
+ N_VSS_c_3_p N_VSS_c_6_p N_VSS_c_9_p N_VSS_c_23_p N_VSS_c_30_p N_VSS_c_10_p
+ N_VSS_c_31_p N_VSS_c_7_p N_VSS_c_8_p N_VSS_c_19_p N_VSS_c_12_p N_VSS_c_20_p
+ N_VSS_c_27_p N_VSS_c_21_p VSS Vss PM_G3_OR2_N1_VSS
x_PM_G3_OR2_N1_VDD N_VDD_XI2.X0_PGD N_VDD_XI2.X0_PGS N_VDD_XI0.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI3.X0_PGD N_VDD_XI3.X0_PGS
+ N_VDD_XI4.X0_S N_VDD_c_78_n N_VDD_c_149_p N_VDD_c_79_n N_VDD_c_140_p
+ N_VDD_c_80_n N_VDD_c_84_n N_VDD_c_88_n N_VDD_c_90_n N_VDD_c_91_n N_VDD_c_124_p
+ N_VDD_c_97_n N_VDD_c_100_n N_VDD_c_104_n N_VDD_c_107_n N_VDD_c_156_p
+ N_VDD_c_112_n N_VDD_c_114_n VDD N_VDD_c_115_n N_VDD_c_116_n N_VDD_c_121_p
+ N_VDD_c_117_n N_VDD_c_119_n Vss PM_G3_OR2_N1_VDD
x_PM_G3_OR2_N1_B N_B_XI2.X0_CG N_B_XI0.X0_CG N_B_c_169_n N_B_c_160_n N_B_c_161_n
+ B N_B_c_164_n N_B_c_165_n Vss PM_G3_OR2_N1_B
x_PM_G3_OR2_N1_NET21 N_NET21_XI2.X0_D N_NET21_XI0.X0_D N_NET21_XI3.X0_CG
+ N_NET21_XI4.X0_CG N_NET21_c_203_n N_NET21_c_190_n N_NET21_c_191_n
+ N_NET21_c_195_n N_NET21_c_212_n N_NET21_c_197_n Vss PM_G3_OR2_N1_NET21
x_PM_G3_OR2_N1_A N_A_XI0.X0_PGS N_A_XI1.X0_CG N_A_c_224_n N_A_c_228_n
+ N_A_c_230_n A Vss PM_G3_OR2_N1_A
x_PM_G3_OR2_N1_Z N_Z_XI3.X0_D Z N_Z_c_248_n Vss PM_G3_OR2_N1_Z
cc_1 N_VSS_XI0.X0_PGD N_VDD_XI1.X0_PGD 0.00175996f
cc_2 N_VSS_XI4.X0_PGD N_VDD_XI3.X0_PGD 0.00168578f
cc_3 N_VSS_c_3_p N_VDD_c_78_n 0.00175996f
cc_4 N_VSS_c_4_p N_VDD_c_79_n 0.00168578f
cc_5 N_VSS_XI2.X0_S N_VDD_c_80_n 9.5668e-19
cc_6 N_VSS_c_6_p N_VDD_c_80_n 0.00165395f
cc_7 N_VSS_c_7_p N_VDD_c_80_n 0.00519974f
cc_8 N_VSS_c_8_p N_VDD_c_80_n 0.00186257f
cc_9 N_VSS_c_9_p N_VDD_c_84_n 4.43871e-19
cc_10 N_VSS_c_10_p N_VDD_c_84_n 3.66936e-19
cc_11 N_VSS_c_7_p N_VDD_c_84_n 0.00303537f
cc_12 N_VSS_c_12_p N_VDD_c_84_n 0.00106607f
cc_13 N_VSS_XI2.X0_S N_VDD_c_88_n 3.7884e-19
cc_14 N_VSS_c_6_p N_VDD_c_88_n 0.00104703f
cc_15 N_VSS_c_6_p N_VDD_c_90_n 7.47067e-19
cc_16 N_VSS_c_3_p N_VDD_c_91_n 3.37151e-19
cc_17 N_VSS_c_9_p N_VDD_c_91_n 0.00161703f
cc_18 N_VSS_c_10_p N_VDD_c_91_n 2.03837e-19
cc_19 N_VSS_c_19_p N_VDD_c_91_n 0.0034844f
cc_20 N_VSS_c_20_p N_VDD_c_91_n 0.00432568f
cc_21 N_VSS_c_21_p N_VDD_c_91_n 7.74609e-19
cc_22 N_VSS_c_9_p N_VDD_c_97_n 8.45115e-19
cc_23 N_VSS_c_23_p N_VDD_c_97_n 3.93845e-19
cc_24 N_VSS_c_10_p N_VDD_c_97_n 3.95933e-19
cc_25 N_VSS_c_23_p N_VDD_c_100_n 5.01863e-19
cc_26 N_VSS_c_20_p N_VDD_c_100_n 0.00137553f
cc_27 N_VSS_c_27_p N_VDD_c_100_n 0.00142235f
cc_28 VSS N_VDD_c_100_n 0.00104966f
cc_29 N_VSS_c_23_p N_VDD_c_104_n 3.91951e-19
cc_30 N_VSS_c_30_p N_VDD_c_104_n 8.51944e-19
cc_31 N_VSS_c_31_p N_VDD_c_104_n 3.99794e-19
cc_32 N_VSS_c_32_p N_VDD_c_107_n 3.80388e-19
cc_33 N_VSS_c_4_p N_VDD_c_107_n 3.60588e-19
cc_34 N_VSS_c_30_p N_VDD_c_107_n 0.00141604f
cc_35 N_VSS_c_31_p N_VDD_c_107_n 0.00112293f
cc_36 N_VSS_c_27_p N_VDD_c_107_n 0.00608608f
cc_37 N_VSS_c_30_p N_VDD_c_112_n 9.12964e-19
cc_38 N_VSS_c_31_p N_VDD_c_112_n 3.66936e-19
cc_39 N_VSS_c_7_p N_VDD_c_114_n 0.00116512f
cc_40 N_VSS_c_20_p N_VDD_c_115_n 9.75006e-19
cc_41 N_VSS_c_27_p N_VDD_c_116_n 9.68945e-19
cc_42 N_VSS_c_9_p N_VDD_c_117_n 3.44698e-19
cc_43 N_VSS_c_10_p N_VDD_c_117_n 7.93802e-19
cc_44 N_VSS_c_30_p N_VDD_c_119_n 3.48267e-19
cc_45 N_VSS_c_31_p N_VDD_c_119_n 8.07896e-19
cc_46 N_VSS_c_10_p N_B_c_160_n 0.00234321f
cc_47 N_VSS_c_9_p N_B_c_161_n 8.39582e-19
cc_48 N_VSS_c_10_p N_B_c_161_n 5.42695e-19
cc_49 N_VSS_c_7_p N_B_c_161_n 7.94601e-19
cc_50 N_VSS_c_10_p N_B_c_164_n 2.00604e-19
cc_51 N_VSS_c_51_p N_B_c_165_n 8.37306e-19
cc_52 N_VSS_c_9_p N_B_c_165_n 4.56568e-19
cc_53 N_VSS_c_10_p N_B_c_165_n 0.00173573f
cc_54 N_VSS_XI2.X0_S N_NET21_XI2.X0_D 3.43419e-19
cc_55 N_VSS_c_6_p N_NET21_XI2.X0_D 3.48267e-19
cc_56 N_VSS_XI1.X0_S N_NET21_XI0.X0_D 3.43419e-19
cc_57 N_VSS_c_23_p N_NET21_XI0.X0_D 3.48267e-19
cc_58 N_VSS_c_31_p N_NET21_XI4.X0_CG 7.99056e-19
cc_59 N_VSS_XI4.X0_PGD N_NET21_c_190_n 4.20799e-19
cc_60 N_VSS_XI1.X0_S N_NET21_c_191_n 3.48267e-19
cc_61 N_VSS_c_6_p N_NET21_c_191_n 8.89782e-19
cc_62 N_VSS_c_23_p N_NET21_c_191_n 5.69026e-19
cc_63 N_VSS_c_7_p N_NET21_c_191_n 2.81358e-19
cc_64 N_VSS_c_7_p N_NET21_c_195_n 2.56803e-19
cc_65 N_VSS_c_27_p N_NET21_c_195_n 2.99166e-19
cc_66 N_VSS_c_23_p N_NET21_c_197_n 9.55513e-19
cc_67 N_VSS_c_7_p N_NET21_c_197_n 2.03357e-19
cc_68 N_VSS_c_20_p N_NET21_c_197_n 9.1856e-19
cc_69 N_VSS_XI0.X0_PGD N_A_c_224_n 9.39677e-19
cc_70 N_VSS_c_3_p N_A_c_224_n 2.16729e-19
cc_71 N_VSS_XI1.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_72 N_VSS_c_23_p N_Z_XI3.X0_D 3.48267e-19
cc_73 N_VSS_XI1.X0_S N_Z_c_248_n 3.48267e-19
cc_74 N_VSS_c_23_p N_Z_c_248_n 7.85754e-19
cc_75 N_VSS_c_27_p N_Z_c_248_n 2.64173e-19
cc_76 N_VDD_c_121_p N_B_XI2.X0_CG 0.00237871f
cc_77 N_VDD_c_121_p N_B_c_169_n 0.00105622f
cc_78 N_VDD_c_80_n N_B_c_161_n 0.0025613f
cc_79 N_VDD_c_124_p N_B_c_161_n 7.31965e-19
cc_80 N_VDD_c_121_p N_B_c_161_n 5.48584e-19
cc_81 N_VDD_c_80_n N_B_c_164_n 4.9897e-19
cc_82 N_VDD_c_124_p N_B_c_164_n 4.85469e-19
cc_83 N_VDD_c_121_p N_B_c_164_n 0.00150793f
cc_84 N_VDD_c_80_n N_B_c_165_n 3.66936e-19
cc_85 N_VDD_c_121_p N_B_c_165_n 2.00604e-19
cc_86 N_VDD_XI0.X0_S N_NET21_XI0.X0_D 3.43419e-19
cc_87 N_VDD_c_90_n N_NET21_XI0.X0_D 3.72199e-19
cc_88 N_VDD_c_91_n N_NET21_XI0.X0_D 3.7884e-19
cc_89 N_VDD_c_119_n N_NET21_c_203_n 0.00250475f
cc_90 N_VDD_XI3.X0_PGD N_NET21_c_190_n 4.25379e-19
cc_91 N_VDD_XI0.X0_S N_NET21_c_191_n 3.48267e-19
cc_92 N_VDD_c_80_n N_NET21_c_191_n 4.38672e-19
cc_93 N_VDD_c_90_n N_NET21_c_191_n 7.89245e-19
cc_94 N_VDD_c_91_n N_NET21_c_191_n 5.36364e-19
cc_95 N_VDD_c_140_p N_NET21_c_195_n 3.64358e-19
cc_96 N_VDD_c_104_n N_NET21_c_195_n 6.84156e-19
cc_97 N_VDD_c_119_n N_NET21_c_195_n 4.99367e-19
cc_98 N_VDD_c_104_n N_NET21_c_212_n 4.85469e-19
cc_99 N_VDD_c_119_n N_NET21_c_212_n 0.0014909f
cc_100 N_VDD_XI2.X0_PGD N_A_c_224_n 5.10213e-19
cc_101 N_VDD_XI1.X0_PGD N_A_c_224_n 2.48727e-19
cc_102 N_VDD_XI2.X0_PGS N_A_c_228_n 6.4837e-19
cc_103 N_VDD_c_80_n N_A_c_228_n 3.16598e-19
cc_104 N_VDD_c_149_p N_A_c_230_n 8.9931e-19
cc_105 N_VDD_c_97_n N_A_c_230_n 4.91217e-19
cc_106 N_VDD_c_117_n N_A_c_230_n 0.00142365f
cc_107 N_VDD_c_97_n A 6.02732e-19
cc_108 N_VDD_c_117_n A 4.56568e-19
cc_109 N_VDD_XI4.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_110 N_VDD_c_107_n N_Z_XI3.X0_D 3.7884e-19
cc_111 N_VDD_c_156_p N_Z_XI3.X0_D 3.72199e-19
cc_112 N_VDD_XI4.X0_S N_Z_c_248_n 3.48267e-19
cc_113 N_VDD_c_107_n N_Z_c_248_n 5.12447e-19
cc_114 N_VDD_c_156_p N_Z_c_248_n 7.4527e-19
cc_115 N_B_c_161_n N_NET21_c_191_n 0.00757794f
cc_116 N_B_c_164_n N_NET21_c_191_n 9.56873e-19
cc_117 N_B_c_165_n N_NET21_c_191_n 8.92526e-19
cc_118 N_B_c_160_n N_A_XI0.X0_PGS 4.5346e-19
cc_119 N_B_c_165_n N_A_XI0.X0_PGS 7.86826e-19
cc_120 N_B_c_164_n N_A_c_224_n 9.25308e-19
cc_121 N_B_c_165_n N_A_c_230_n 7.50183e-19
cc_122 N_NET21_c_191_n N_A_c_224_n 8.63036e-19
cc_123 N_NET21_c_191_n N_A_c_230_n 9.38449e-19
cc_124 N_NET21_c_195_n N_A_c_230_n 3.48267e-19
cc_125 N_NET21_c_212_n N_A_c_230_n 0.00196751f
cc_126 N_NET21_c_191_n A 0.00142917f
cc_127 N_NET21_c_195_n A 4.28721e-19
cc_128 N_NET21_c_197_n A 3.26205e-19
*
.ends
*
*
.subckt OR2_HPNW4 A B Y VDD VSS
xgate (VSS VDD B A Y) G3_OR2_N1_2
.ends
*
* File: G4_XNOR2_N1.pex.netlist
* Created: Wed Mar 16 10:29:55 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*







.subckt G4_XNOR2_N1_2 VDD VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI1.X0 N_NET1_XI1.X0_D N_VSS_XI1.X0_PGD N_B_XI1.X0_CG N_VSS_XI1.X0_PGD
+ N_VDD_XI1.X0_S TIGFET_HPNW4
XI9.X0 N_NET2_XI9.X0_D N_VDD_XI9.X0_PGD N_A_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI10.X0 N_NET1_XI1.X0_D N_VDD_XI10.X0_PGD N_B_XI10.X0_CG N_VDD_XI10.X0_PGD
+ N_VSS_XI10.X0_S TIGFET_HPNW4
XI3.X0 N_NET2_XI9.X0_D N_VSS_XI3.X0_PGD N_A_XI3.X0_CG N_VSS_XI3.X0_PGD
+ N_VDD_XI3.X0_S TIGFET_HPNW4
XI5.X0 N_Z_XI5.X0_D N_B_XI5.X0_PGD N_NET2_XI5.X0_CG N_B_XI5.X0_PGD
+ N_VSS_XI10.X0_S TIGFET_HPNW4
XI8.X0 N_Z_XI8.X0_D N_A_XI8.X0_PGD N_B_XI8.X0_CG N_A_XI8.X0_PGD N_VDD_XI3.X0_S
+ TIGFET_HPNW4
XI11.X0 N_Z_XI5.X0_D N_NET1_XI11.X0_PGD N_A_XI11.X0_CG N_NET1_XI11.X0_PGD
+ N_VSS_XI11.X0_S TIGFET_HPNW4
XI7.X0 N_Z_XI8.X0_D N_NET2_XI7.X0_PGD N_NET1_XI7.X0_CG N_NET2_XI7.X0_PGD
+ N_VDD_XI7.X0_S TIGFET_HPNW4
*
x_PM_G4_XNOR2_N1_VDD N_VDD_XI1.X0_S N_VDD_XI9.X0_PGD N_VDD_XI10.X0_PGD
+ N_VDD_XI3.X0_S N_VDD_XI7.X0_S N_VDD_c_11_p N_VDD_c_58_p N_VDD_c_26_p
+ N_VDD_c_8_p N_VDD_c_17_p N_VDD_c_14_p N_VDD_c_9_p N_VDD_c_45_p N_VDD_c_3_p
+ N_VDD_c_16_p N_VDD_c_49_p N_VDD_c_21_p N_VDD_c_12_p N_VDD_c_19_p N_VDD_c_4_p
+ N_VDD_c_60_p N_VDD_c_7_p N_VDD_c_90_p N_VDD_c_42_p N_VDD_c_48_p VDD
+ N_VDD_c_24_p N_VDD_c_20_p Vss PM_G4_XNOR2_N1_VDD
x_PM_G4_XNOR2_N1_VSS N_VSS_XI1.X0_PGD N_VSS_XI9.X0_S N_VSS_XI10.X0_S
+ N_VSS_XI3.X0_PGD N_VSS_XI11.X0_S N_VSS_c_121_n N_VSS_c_123_n N_VSS_c_172_p
+ N_VSS_c_124_n N_VSS_c_126_n N_VSS_c_130_n N_VSS_c_134_n N_VSS_c_138_n
+ N_VSS_c_143_n N_VSS_c_145_n N_VSS_c_149_n N_VSS_c_153_n N_VSS_c_156_n
+ N_VSS_c_157_n N_VSS_c_158_n N_VSS_c_159_n N_VSS_c_162_n N_VSS_c_163_n
+ N_VSS_c_164_n N_VSS_c_185_p N_VSS_c_165_n N_VSS_c_166_n VSS Vss
+ PM_G4_XNOR2_N1_VSS
x_PM_G4_XNOR2_N1_A N_A_XI9.X0_CG N_A_XI3.X0_CG N_A_XI8.X0_PGD N_A_XI11.X0_CG
+ N_A_c_214_n N_A_c_215_n N_A_c_217_n N_A_c_218_n N_A_c_249_p N_A_c_219_n
+ N_A_c_220_n A N_A_c_223_n N_A_c_225_n N_A_c_226_n N_A_c_229_n N_A_c_244_p
+ N_A_c_242_n Vss PM_G4_XNOR2_N1_A
x_PM_G4_XNOR2_N1_NET1 N_NET1_XI1.X0_D N_NET1_XI11.X0_PGD N_NET1_XI7.X0_CG
+ N_NET1_c_309_p N_NET1_c_293_n N_NET1_c_276_n N_NET1_c_279_n N_NET1_c_296_n
+ N_NET1_c_280_n Vss PM_G4_XNOR2_N1_NET1
x_PM_G4_XNOR2_N1_NET2 N_NET2_XI9.X0_D N_NET2_XI5.X0_CG N_NET2_XI7.X0_PGD
+ N_NET2_c_336_n N_NET2_c_356_p N_NET2_c_314_n N_NET2_c_315_n N_NET2_c_318_n
+ N_NET2_c_322_n N_NET2_c_324_n Vss PM_G4_XNOR2_N1_NET2
x_PM_G4_XNOR2_N1_B N_B_XI1.X0_CG N_B_XI10.X0_CG N_B_XI5.X0_PGD N_B_XI8.X0_CG
+ N_B_c_363_n N_B_c_382_n N_B_c_365_n N_B_c_392_n N_B_c_388_n N_B_c_384_n
+ N_B_c_395_n N_B_c_366_n N_B_c_367_n B N_B_c_369_n Vss PM_G4_XNOR2_N1_B
x_PM_G4_XNOR2_N1_Z N_Z_XI5.X0_D N_Z_XI8.X0_D N_Z_c_403_n Z Vss PM_G4_XNOR2_N1_Z
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI1.X0_PGD 2.96813e-19
cc_2 N_VDD_XI10.X0_PGD N_VSS_XI1.X0_PGD 0.00168295f
cc_3 N_VDD_c_3_p N_VSS_XI9.X0_S 2.15082e-19
cc_4 N_VDD_c_4_p N_VSS_XI10.X0_S 2.35318e-19
cc_5 N_VDD_XI9.X0_PGD N_VSS_XI3.X0_PGD 0.00167677f
cc_6 N_VDD_c_4_p N_VSS_XI3.X0_PGD 2.68479e-19
cc_7 N_VDD_c_7_p N_VSS_XI11.X0_S 2.15082e-19
cc_8 N_VDD_c_8_p N_VSS_c_121_n 0.00168295f
cc_9 N_VDD_c_9_p N_VSS_c_121_n 3.60588e-19
cc_10 N_VDD_c_9_p N_VSS_c_123_n 3.60588e-19
cc_11 N_VDD_c_11_p N_VSS_c_124_n 0.00167677f
cc_12 N_VDD_c_12_p N_VSS_c_124_n 3.60588e-19
cc_13 N_VDD_XI1.X0_S N_VSS_c_126_n 2.15082e-19
cc_14 N_VDD_c_14_p N_VSS_c_126_n 0.00187494f
cc_15 N_VDD_c_3_p N_VSS_c_126_n 8.9077e-19
cc_16 N_VDD_c_16_p N_VSS_c_126_n 5.16845e-19
cc_17 N_VDD_c_17_p N_VSS_c_130_n 4.43871e-19
cc_18 N_VDD_c_9_p N_VSS_c_130_n 0.00141228f
cc_19 N_VDD_c_19_p N_VSS_c_130_n 8.52111e-19
cc_20 N_VDD_c_20_p N_VSS_c_130_n 3.48267e-19
cc_21 N_VDD_c_21_p N_VSS_c_134_n 9.21268e-19
cc_22 N_VDD_c_12_p N_VSS_c_134_n 0.00141228f
cc_23 N_VDD_c_4_p N_VSS_c_134_n 0.00225084f
cc_24 N_VDD_c_24_p N_VSS_c_134_n 3.48267e-19
cc_25 N_VDD_XI3.X0_S N_VSS_c_138_n 2.35318e-19
cc_26 N_VDD_c_26_p N_VSS_c_138_n 2.72094e-19
cc_27 N_VDD_c_9_p N_VSS_c_138_n 0.00534617f
cc_28 N_VDD_c_4_p N_VSS_c_138_n 4.25159e-19
cc_29 N_VDD_c_20_p N_VSS_c_138_n 9.58524e-19
cc_30 N_VDD_XI7.X0_S N_VSS_c_143_n 2.15082e-19
cc_31 N_VDD_c_7_p N_VSS_c_143_n 3.16299e-19
cc_32 N_VDD_c_17_p N_VSS_c_145_n 3.66936e-19
cc_33 N_VDD_c_9_p N_VSS_c_145_n 0.00112249f
cc_34 N_VDD_c_19_p N_VSS_c_145_n 3.99794e-19
cc_35 N_VDD_c_20_p N_VSS_c_145_n 8.03027e-19
cc_36 N_VDD_c_21_p N_VSS_c_149_n 3.82294e-19
cc_37 N_VDD_c_12_p N_VSS_c_149_n 0.00112249f
cc_38 N_VDD_c_4_p N_VSS_c_149_n 9.55322e-19
cc_39 N_VDD_c_24_p N_VSS_c_149_n 8.0279e-19
cc_40 N_VDD_c_17_p N_VSS_c_153_n 0.00287902f
cc_41 N_VDD_c_14_p N_VSS_c_153_n 0.0057117f
cc_42 N_VDD_c_42_p N_VSS_c_153_n 0.0010706f
cc_43 N_VDD_c_14_p N_VSS_c_156_n 0.00304013f
cc_44 N_VDD_c_9_p N_VSS_c_157_n 0.00342836f
cc_45 N_VDD_c_45_p N_VSS_c_158_n 0.00107429f
cc_46 N_VDD_c_16_p N_VSS_c_159_n 0.00352516f
cc_47 N_VDD_c_12_p N_VSS_c_159_n 0.0060405f
cc_48 N_VDD_c_48_p N_VSS_c_159_n 0.00101104f
cc_49 N_VDD_c_49_p N_VSS_c_162_n 0.00105833f
cc_50 N_VDD_c_9_p N_VSS_c_163_n 0.00458401f
cc_51 N_VDD_c_7_p N_VSS_c_164_n 0.00135143f
cc_52 N_VDD_c_14_p N_VSS_c_165_n 7.88896e-19
cc_53 N_VDD_c_9_p N_VSS_c_166_n 7.74609e-19
cc_54 N_VDD_c_4_p N_A_XI8.X0_PGD 2.51969e-19
cc_55 N_VDD_c_24_p N_A_c_214_n 0.00237738f
cc_56 N_VDD_XI9.X0_PGD N_A_c_215_n 4.04053e-19
cc_57 N_VDD_XI10.X0_PGD N_A_c_215_n 2.40582e-19
cc_58 N_VDD_c_58_p N_A_c_217_n 9.54306e-19
cc_59 N_VDD_XI10.X0_PGD N_A_c_218_n 2.40582e-19
cc_60 N_VDD_c_60_p N_A_c_219_n 5.838e-19
cc_61 N_VDD_c_14_p N_A_c_220_n 5.24876e-19
cc_62 N_VDD_c_21_p N_A_c_220_n 6.41525e-19
cc_63 N_VDD_c_24_p N_A_c_220_n 4.56568e-19
cc_64 N_VDD_c_4_p N_A_c_223_n 0.00237851f
cc_65 N_VDD_c_60_p N_A_c_223_n 0.00200281f
cc_66 N_VDD_c_60_p N_A_c_225_n 8.17097e-19
cc_67 N_VDD_c_14_p N_A_c_226_n 6.27972e-19
cc_68 N_VDD_c_21_p N_A_c_226_n 4.85469e-19
cc_69 N_VDD_c_24_p N_A_c_226_n 6.1245e-19
cc_70 N_VDD_c_4_p N_A_c_229_n 9.84209e-19
cc_71 N_VDD_c_60_p N_A_c_229_n 2.37583e-19
cc_72 N_VDD_XI1.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_73 N_VDD_c_9_p N_NET1_XI1.X0_D 3.7884e-19
cc_74 N_VDD_c_3_p N_NET1_XI1.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_S N_NET1_c_276_n 3.48267e-19
cc_76 N_VDD_c_9_p N_NET1_c_276_n 4.58491e-19
cc_77 N_VDD_c_3_p N_NET1_c_276_n 5.226e-19
cc_78 N_VDD_c_19_p N_NET1_c_279_n 0.00121121f
cc_79 N_VDD_c_9_p N_NET1_c_280_n 3.78572e-19
cc_80 N_VDD_XI3.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_81 N_VDD_c_12_p N_NET2_XI9.X0_D 3.7884e-19
cc_82 N_VDD_c_4_p N_NET2_XI9.X0_D 3.48267e-19
cc_83 N_VDD_c_60_p N_NET2_c_314_n 8.01015e-19
cc_84 N_VDD_XI3.X0_S N_NET2_c_315_n 3.48267e-19
cc_85 N_VDD_c_12_p N_NET2_c_315_n 4.58491e-19
cc_86 N_VDD_c_4_p N_NET2_c_315_n 8.45449e-19
cc_87 N_VDD_c_12_p N_NET2_c_318_n 3.29894e-19
cc_88 N_VDD_c_4_p N_NET2_c_318_n 8.51778e-19
cc_89 N_VDD_c_60_p N_NET2_c_318_n 0.00334727f
cc_90 N_VDD_c_90_p N_NET2_c_318_n 7.7731e-19
cc_91 N_VDD_c_60_p N_NET2_c_322_n 2.33029e-19
cc_92 N_VDD_c_90_p N_NET2_c_322_n 3.66936e-19
cc_93 N_VDD_c_21_p N_NET2_c_324_n 3.10284e-19
cc_94 N_VDD_c_20_p N_B_XI10.X0_CG 0.00237871f
cc_95 N_VDD_XI10.X0_PGD N_B_XI5.X0_PGD 0.00176522f
cc_96 N_VDD_XI9.X0_PGD N_B_c_363_n 2.40582e-19
cc_97 N_VDD_XI10.X0_PGD N_B_c_363_n 4.04053e-19
cc_98 N_VDD_XI10.X0_PGD N_B_c_365_n 4.05198e-19
cc_99 N_VDD_c_26_p N_B_c_366_n 0.00154836f
cc_100 N_VDD_c_19_p N_B_c_367_n 5.50671e-19
cc_101 N_VDD_c_20_p N_B_c_367_n 8.9014e-19
cc_102 N_VDD_c_19_p N_B_c_369_n 4.73723e-19
cc_103 N_VDD_c_20_p N_B_c_369_n 0.0014909f
cc_104 N_VDD_XI3.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_105 N_VDD_XI7.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_106 N_VDD_c_4_p N_Z_XI8.X0_D 3.48267e-19
cc_107 N_VDD_c_60_p N_Z_XI8.X0_D 3.7884e-19
cc_108 N_VDD_c_7_p N_Z_XI8.X0_D 3.72199e-19
cc_109 N_VDD_XI3.X0_S N_Z_c_403_n 3.48267e-19
cc_110 N_VDD_XI7.X0_S N_Z_c_403_n 3.48267e-19
cc_111 N_VDD_c_4_p N_Z_c_403_n 5.21254e-19
cc_112 N_VDD_c_60_p N_Z_c_403_n 6.55718e-19
cc_113 N_VDD_c_7_p N_Z_c_403_n 8.25922e-19
cc_114 N_VSS_c_149_n N_A_XI3.X0_CG 9.02944e-19
cc_115 N_VSS_XI3.X0_PGD N_A_XI8.X0_PGD 0.00150976f
cc_116 N_VSS_XI1.X0_PGD N_A_c_215_n 2.40582e-19
cc_117 N_VSS_XI3.X0_PGD N_A_c_215_n 3.99472e-19
cc_118 N_VSS_XI3.X0_PGD N_A_c_218_n 4.05198e-19
cc_119 N_VSS_c_172_p N_A_c_219_n 0.00150976f
cc_120 N_VSS_c_134_n N_A_c_223_n 4.12959e-19
cc_121 N_VSS_c_153_n N_A_c_223_n 3.96361e-19
cc_122 N_VSS_c_163_n N_A_c_225_n 2.41875e-19
cc_123 N_VSS_c_145_n N_A_c_226_n 4.65658e-19
cc_124 N_VSS_c_149_n N_A_c_229_n 8.90609e-19
cc_125 N_VSS_c_163_n N_A_c_242_n 3.10545e-19
cc_126 N_VSS_XI10.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_127 N_VSS_c_138_n N_NET1_XI1.X0_D 3.48267e-19
cc_128 N_VSS_XI10.X0_S N_NET1_c_276_n 3.48267e-19
cc_129 N_VSS_c_138_n N_NET1_c_276_n 0.0012813f
cc_130 N_VSS_c_138_n N_NET1_c_279_n 0.00174104f
cc_131 N_VSS_c_163_n N_NET1_c_279_n 5.89244e-19
cc_132 N_VSS_c_185_p N_NET1_c_279_n 0.00121599f
cc_133 N_VSS_c_130_n N_NET1_c_280_n 0.00206231f
cc_134 N_VSS_c_153_n N_NET1_c_280_n 9.32604e-19
cc_135 N_VSS_c_163_n N_NET1_c_280_n 0.0214545f
cc_136 N_VSS_XI9.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_137 N_VSS_c_126_n N_NET2_XI9.X0_D 3.48267e-19
cc_138 N_VSS_XI9.X0_S N_NET2_c_315_n 3.48267e-19
cc_139 N_VSS_c_126_n N_NET2_c_315_n 0.00108327f
cc_140 N_VSS_c_159_n N_NET2_c_315_n 3.31434e-19
cc_141 N_VSS_c_134_n N_NET2_c_318_n 0.00143089f
cc_142 N_VSS_c_156_n N_NET2_c_324_n 3.36104e-19
cc_143 N_VSS_c_159_n N_NET2_c_324_n 6.48614e-19
cc_144 N_VSS_c_145_n N_B_XI1.X0_CG 9.02944e-19
cc_145 N_VSS_XI1.X0_PGD N_B_c_363_n 3.99472e-19
cc_146 N_VSS_XI3.X0_PGD N_B_c_363_n 2.40582e-19
cc_147 N_VSS_XI3.X0_PGD N_B_c_365_n 2.40582e-19
cc_148 N_VSS_c_138_n N_B_c_366_n 2.8419e-19
cc_149 N_VSS_c_149_n N_B_c_367_n 2.07877e-19
cc_150 N_VSS_c_153_n N_B_c_367_n 2.27769e-19
cc_151 N_VSS_c_149_n N_B_c_369_n 7.33679e-19
cc_152 N_VSS_XI10.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_153 N_VSS_XI11.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_154 N_VSS_c_138_n N_Z_XI5.X0_D 3.48267e-19
cc_155 N_VSS_c_143_n N_Z_XI5.X0_D 3.48267e-19
cc_156 N_VSS_XI10.X0_S N_Z_c_403_n 3.48267e-19
cc_157 N_VSS_XI11.X0_S N_Z_c_403_n 3.48267e-19
cc_158 N_VSS_c_138_n N_Z_c_403_n 8.61925e-19
cc_159 N_VSS_c_143_n N_Z_c_403_n 5.69026e-19
cc_160 N_A_XI11.X0_CG N_NET1_XI11.X0_PGD 4.5346e-19
cc_161 N_A_c_244_p N_NET1_XI11.X0_PGD 0.00151381f
cc_162 N_A_c_244_p N_NET1_c_293_n 0.00157635f
cc_163 N_A_c_225_n N_NET1_c_279_n 0.00310276f
cc_164 N_A_c_242_n N_NET1_c_279_n 0.00205512f
cc_165 N_A_XI11.X0_CG N_NET1_c_296_n 0.00234108f
cc_166 N_A_c_249_p N_NET1_c_296_n 0.00101616f
cc_167 N_A_c_244_p N_NET1_c_296_n 0.00161406f
cc_168 N_A_XI8.X0_PGD N_NET2_XI7.X0_PGD 0.00160287f
cc_169 N_A_c_218_n N_NET2_XI7.X0_PGD 3.14428e-19
cc_170 N_A_c_244_p N_NET2_XI7.X0_PGD 5.68075e-19
cc_171 N_A_XI8.X0_PGD N_NET2_c_336_n 4.60549e-19
cc_172 N_A_c_219_n N_NET2_c_314_n 0.00160287f
cc_173 N_A_c_223_n N_NET2_c_315_n 7.37727e-19
cc_174 N_A_c_223_n N_NET2_c_318_n 0.00205074f
cc_175 N_A_c_225_n N_NET2_c_318_n 0.0018485f
cc_176 N_A_c_229_n N_NET2_c_318_n 3.44698e-19
cc_177 N_A_c_223_n N_NET2_c_322_n 3.44698e-19
cc_178 N_A_c_229_n N_NET2_c_322_n 9.07485e-19
cc_179 N_A_c_244_p N_NET2_c_322_n 3.98239e-19
cc_180 N_A_c_218_n N_B_XI8.X0_CG 0.003858f
cc_181 N_A_c_229_n N_B_XI8.X0_CG 0.00111269f
cc_182 N_A_c_215_n N_B_c_363_n 0.00575421f
cc_183 N_A_c_226_n N_B_c_382_n 4.09767e-19
cc_184 N_A_c_218_n N_B_c_365_n 0.00308843f
cc_185 N_A_c_218_n N_B_c_384_n 0.00362155f
cc_186 N_A_c_215_n N_B_c_369_n 6.77269e-19
cc_187 N_A_c_223_n N_Z_c_403_n 0.00321233f
cc_188 N_A_c_225_n N_Z_c_403_n 0.0025035f
cc_189 N_A_c_244_p N_Z_c_403_n 8.50872e-19
cc_190 N_NET1_c_276_n N_NET2_XI9.X0_D 2.15082e-19
cc_191 N_NET1_XI11.X0_PGD N_NET2_XI5.X0_CG 2.62058e-19
cc_192 N_NET1_c_293_n N_NET2_XI7.X0_PGD 0.00832016f
cc_193 N_NET1_XI11.X0_PGD N_NET2_c_336_n 0.00416722f
cc_194 N_NET1_XI1.X0_D N_NET2_c_315_n 2.15082e-19
cc_195 N_NET1_c_279_n N_NET2_c_318_n 0.00142494f
cc_196 N_NET1_XI7.X0_CG N_NET2_c_322_n 0.00102831f
cc_197 N_NET1_XI11.X0_PGD N_B_XI5.X0_PGD 0.00188492f
cc_198 N_NET1_XI7.X0_CG N_B_XI8.X0_CG 2.60667e-19
cc_199 N_NET1_c_293_n N_B_c_388_n 2.60667e-19
cc_200 N_NET1_c_309_p N_B_c_366_n 0.00165894f
cc_201 N_NET1_c_279_n N_Z_c_403_n 3.02205e-19
cc_202 N_NET2_XI5.X0_CG N_B_XI5.X0_PGD 0.0019183f
cc_203 N_NET2_c_336_n N_B_XI5.X0_PGD 0.00161994f
cc_204 N_NET2_XI7.X0_PGD N_B_c_392_n 3.1641e-19
cc_205 N_NET2_XI7.X0_PGD N_B_c_388_n 0.00313953f
cc_206 N_NET2_c_356_p N_B_c_388_n 0.00172424f
cc_207 N_NET2_c_356_p N_B_c_395_n 0.0019183f
cc_208 N_NET2_XI7.X0_PGD N_Z_c_403_n 0.00115814f
cc_209 N_NET2_c_336_n N_Z_c_403_n 5.21666e-19
cc_210 N_NET2_c_318_n N_Z_c_403_n 2.80086e-19
cc_211 N_B_c_388_n N_Z_c_403_n 8.84927e-19
cc_212 N_B_c_367_n N_Z_c_403_n 3.17615e-19
*
.ends
*
*
.subckt XNOR2_HPNW4 A B Y VDD VSS
xgate (VDD VSS A B Y) G4_XNOR2_N1_2
.ends
*
* File: G5_XNOR3_N1.pex.netlist
* Created: Fri Mar 25 15:42:00 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*









.subckt G5_XNOR3_N1_2 VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI10.X0 N_CI_XI10.X0_D N_VSS_XI10.X0_PGD N_C_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW4
XI9.X0 N_CI_XI10.X0_D N_VDD_XI9.X0_PGD N_C_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI5.X0 N_BI_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI6.X0 N_BI_XI5.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW4
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW4
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_B_XI2.X0_CG N_AI_XI2.X0_PGD N_C_XI2.X0_S
+ TIGFET_HPNW4
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_BI_XI4.X0_CG N_AI_XI4.X0_PGD N_CI_XI4.X0_S
+ TIGFET_HPNW4
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_BI_XI3.X0_CG N_A_XI3.X0_PGD N_C_XI3.X0_S
+ TIGFET_HPNW4
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_B_XI1.X0_CG N_A_XI1.X0_PGD N_CI_XI1.X0_S
+ TIGFET_HPNW4
*
x_PM_G5_XNOR3_N1_VDD N_VDD_XI10.X0_S N_VDD_XI9.X0_PGD N_VDD_XI5.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI6.X0_S N_VDD_XI7.X0_PGD N_VDD_c_120_p N_VDD_c_18_p
+ N_VDD_c_23_p N_VDD_c_4_p N_VDD_c_110_p N_VDD_c_19_p N_VDD_c_6_p N_VDD_c_25_p
+ N_VDD_c_5_p N_VDD_c_64_p N_VDD_c_27_p N_VDD_c_28_p N_VDD_c_29_p N_VDD_c_35_p
+ N_VDD_c_32_p N_VDD_c_20_p N_VDD_c_11_p N_VDD_c_24_p N_VDD_c_37_p N_VDD_c_12_p
+ N_VDD_c_60_p VDD N_VDD_c_68_p N_VDD_c_72_p N_VDD_c_2_p N_VDD_c_42_p
+ N_VDD_c_38_p Vss PM_G5_XNOR3_N1_VDD
x_PM_G5_XNOR3_N1_C N_C_XI10.X0_CG N_C_XI9.X0_CG N_C_XI2.X0_S N_C_XI3.X0_S
+ N_C_c_143_p N_C_c_125_n N_C_c_136_p C N_C_c_138_p N_C_c_158_p N_C_c_178_p
+ N_C_c_130_n N_C_c_132_n N_C_c_133_n N_C_c_156_p N_C_c_139_p N_C_c_161_p Vss
+ PM_G5_XNOR3_N1_C
x_PM_G5_XNOR3_N1_VSS N_VSS_XI10.X0_PGD N_VSS_XI9.X0_S N_VSS_XI8.X0_PGD
+ N_VSS_XI6.X0_PGD N_VSS_XI7.X0_S N_VSS_c_188_n N_VSS_c_247_n N_VSS_c_189_n
+ N_VSS_c_191_n N_VSS_c_287_p N_VSS_c_192_n N_VSS_c_193_n N_VSS_c_195_n
+ N_VSS_c_201_n N_VSS_c_205_n N_VSS_c_209_n N_VSS_c_213_n N_VSS_c_216_n
+ N_VSS_c_217_n N_VSS_c_220_n N_VSS_c_224_n N_VSS_c_228_n N_VSS_c_231_n
+ N_VSS_c_233_n N_VSS_c_234_n N_VSS_c_235_n N_VSS_c_239_n N_VSS_c_240_n VSS
+ N_VSS_c_243_n N_VSS_c_244_n N_VSS_c_245_n Vss PM_G5_XNOR3_N1_VSS
x_PM_G5_XNOR3_N1_CI N_CI_XI10.X0_D N_CI_XI4.X0_S N_CI_XI1.X0_S N_CI_c_316_n
+ N_CI_c_334_n N_CI_c_356_p N_CI_c_320_n N_CI_c_338_n N_CI_c_324_n N_CI_c_349_p
+ Vss PM_G5_XNOR3_N1_CI
x_PM_G5_XNOR3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI3.X0_PGD N_A_XI1.X0_PGD
+ N_A_c_387_n N_A_c_362_n N_A_c_415_p N_A_c_417_p N_A_c_363_n A N_A_c_370_n
+ N_A_c_381_n N_A_c_371_n N_A_c_372_n N_A_c_386_n N_A_c_374_n N_A_c_399_p Vss
+ PM_G5_XNOR3_N1_A
x_PM_G5_XNOR3_N1_BI N_BI_XI5.X0_D N_BI_XI4.X0_CG N_BI_XI3.X0_CG N_BI_c_478_p
+ N_BI_c_465_n N_BI_c_443_n N_BI_c_468_n N_BI_c_459_n N_BI_c_471_n N_BI_c_472_n
+ N_BI_c_447_n N_BI_c_457_n N_BI_c_477_n N_BI_c_450_n N_BI_c_503_p N_BI_c_451_n
+ Vss PM_G5_XNOR3_N1_BI
x_PM_G5_XNOR3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_523_n
+ N_AI_c_546_n N_AI_c_513_n N_AI_c_514_n N_AI_c_517_n N_AI_c_528_n N_AI_c_518_n
+ Vss PM_G5_XNOR3_N1_AI
x_PM_G5_XNOR3_N1_B N_B_XI5.X0_CG N_B_XI6.X0_CG N_B_XI2.X0_CG N_B_XI1.X0_CG
+ N_B_c_559_n N_B_c_561_n N_B_c_571_n N_B_c_580_n N_B_c_581_n B N_B_c_584_n
+ N_B_c_575_n N_B_c_562_n N_B_c_589_n N_B_c_590_n N_B_c_563_n N_B_c_607_n
+ N_B_c_576_n Vss PM_G5_XNOR3_N1_B
x_PM_G5_XNOR3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_624_n Z Vss PM_G5_XNOR3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_C_XI9.X0_CG 9.58934e-19
cc_2 N_VDD_c_2_p N_C_XI9.X0_CG 8.03148e-19
cc_3 N_VDD_XI9.X0_PGD N_C_c_125_n 4.16623e-19
cc_4 N_VDD_c_4_p N_C_c_125_n 9.58934e-19
cc_5 N_VDD_c_5_p N_C_c_125_n 0.00125128f
cc_6 N_VDD_c_6_p C 3.00172e-19
cc_7 N_VDD_c_5_p C 0.00118142f
cc_8 N_VDD_c_6_p N_C_c_130_n 4.71537e-19
cc_9 N_VDD_c_5_p N_C_c_130_n 2.74773e-19
cc_10 N_VDD_XI6.X0_S N_C_c_132_n 3.43419e-19
cc_11 N_VDD_c_11_p N_C_c_133_n 5.30636e-19
cc_12 N_VDD_c_12_p N_C_c_133_n 7.99481e-19
cc_13 N_VDD_XI9.X0_PGD N_VSS_XI10.X0_PGD 0.00173038f
cc_14 N_VDD_XI5.X0_PGD N_VSS_XI8.X0_PGD 2.27468e-19
cc_15 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172039f
cc_16 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017188f
cc_17 N_VDD_XI7.X0_PGD N_VSS_XI6.X0_PGD 2.1536e-19
cc_18 N_VDD_c_18_p N_VSS_c_188_n 0.00173038f
cc_19 N_VDD_c_19_p N_VSS_c_189_n 0.00172039f
cc_20 N_VDD_c_20_p N_VSS_c_189_n 2.46461e-19
cc_21 N_VDD_c_20_p N_VSS_c_191_n 3.60588e-19
cc_22 N_VDD_c_12_p N_VSS_c_192_n 2.35445e-19
cc_23 N_VDD_c_23_p N_VSS_c_193_n 0.0017188f
cc_24 N_VDD_c_24_p N_VSS_c_193_n 2.74208e-19
cc_25 N_VDD_c_25_p N_VSS_c_195_n 4.32468e-19
cc_26 N_VDD_c_5_p N_VSS_c_195_n 4.60511e-19
cc_27 N_VDD_c_27_p N_VSS_c_195_n 0.00130521f
cc_28 N_VDD_c_28_p N_VSS_c_195_n 4.50568e-19
cc_29 N_VDD_c_29_p N_VSS_c_195_n 3.98949e-19
cc_30 N_VDD_c_2_p N_VSS_c_195_n 3.48267e-19
cc_31 N_VDD_c_5_p N_VSS_c_201_n 5.01863e-19
cc_32 N_VDD_c_32_p N_VSS_c_201_n 2.14355e-19
cc_33 N_VDD_c_11_p N_VSS_c_201_n 7.9087e-19
cc_34 N_VDD_c_12_p N_VSS_c_201_n 3.30117e-19
cc_35 N_VDD_c_35_p N_VSS_c_205_n 6.99368e-19
cc_36 N_VDD_c_20_p N_VSS_c_205_n 0.00161703f
cc_37 N_VDD_c_37_p N_VSS_c_205_n 8.32098e-19
cc_38 N_VDD_c_38_p N_VSS_c_205_n 3.48267e-19
cc_39 N_VDD_c_11_p N_VSS_c_209_n 6.79271e-19
cc_40 N_VDD_c_24_p N_VSS_c_209_n 0.00161703f
cc_41 N_VDD_c_12_p N_VSS_c_209_n 0.00241473f
cc_42 N_VDD_c_42_p N_VSS_c_209_n 3.48267e-19
cc_43 N_VDD_XI7.X0_PGD N_VSS_c_213_n 3.41313e-19
cc_44 N_VDD_c_37_p N_VSS_c_213_n 0.00506009f
cc_45 N_VDD_c_38_p N_VSS_c_213_n 9.58524e-19
cc_46 N_VDD_c_20_p N_VSS_c_216_n 0.00415364f
cc_47 N_VDD_c_25_p N_VSS_c_217_n 4.41003e-19
cc_48 N_VDD_c_29_p N_VSS_c_217_n 3.89161e-19
cc_49 N_VDD_c_2_p N_VSS_c_217_n 7.99831e-19
cc_50 N_VDD_c_35_p N_VSS_c_220_n 3.48267e-19
cc_51 N_VDD_c_20_p N_VSS_c_220_n 2.03837e-19
cc_52 N_VDD_c_37_p N_VSS_c_220_n 3.99794e-19
cc_53 N_VDD_c_38_p N_VSS_c_220_n 8.03027e-19
cc_54 N_VDD_c_11_p N_VSS_c_224_n 3.82294e-19
cc_55 N_VDD_c_24_p N_VSS_c_224_n 2.03837e-19
cc_56 N_VDD_c_12_p N_VSS_c_224_n 9.55109e-19
cc_57 N_VDD_c_42_p N_VSS_c_224_n 8.01441e-19
cc_58 N_VDD_c_6_p N_VSS_c_228_n 0.00301593f
cc_59 N_VDD_c_25_p N_VSS_c_228_n 7.60301e-19
cc_60 N_VDD_c_60_p N_VSS_c_228_n 0.0010705f
cc_61 N_VDD_c_25_p N_VSS_c_231_n 0.00803422f
cc_62 N_VDD_c_29_p N_VSS_c_231_n 8.94414e-19
cc_63 N_VDD_c_5_p N_VSS_c_233_n 0.00969041f
cc_64 N_VDD_c_64_p N_VSS_c_234_n 0.00107143f
cc_65 N_VDD_c_28_p N_VSS_c_235_n 0.00807788f
cc_66 N_VDD_c_32_p N_VSS_c_235_n 7.22996e-19
cc_67 N_VDD_c_20_p N_VSS_c_235_n 0.00374557f
cc_68 N_VDD_c_68_p N_VSS_c_235_n 0.00137227f
cc_69 N_VDD_c_25_p N_VSS_c_239_n 0.00107355f
cc_70 N_VDD_c_5_p N_VSS_c_240_n 0.00142851f
cc_71 N_VDD_c_24_p N_VSS_c_240_n 0.00577339f
cc_72 N_VDD_c_72_p N_VSS_c_240_n 0.00106333f
cc_73 N_VDD_c_25_p N_VSS_c_243_n 0.00112682f
cc_74 N_VDD_c_5_p N_VSS_c_244_n 0.00104966f
cc_75 N_VDD_c_20_p N_VSS_c_245_n 7.74609e-19
cc_76 N_VDD_XI10.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_77 N_VDD_c_27_p N_CI_XI10.X0_D 3.72199e-19
cc_78 N_VDD_XI10.X0_S N_CI_c_316_n 3.48267e-19
cc_79 N_VDD_c_5_p N_CI_c_316_n 5.01863e-19
cc_80 N_VDD_c_27_p N_CI_c_316_n 5.226e-19
cc_81 N_VDD_c_29_p N_CI_c_316_n 0.00213742f
cc_82 N_VDD_c_35_p N_CI_c_320_n 7.47076e-19
cc_83 N_VDD_c_32_p N_CI_c_320_n 4.06004e-19
cc_84 N_VDD_c_38_p N_A_XI7.X0_CG 9.92565e-19
cc_85 N_VDD_XI7.X0_PGD N_A_c_362_n 3.90792e-19
cc_86 N_VDD_XI6.X0_S N_A_c_363_n 2.96819e-19
cc_87 N_VDD_XI7.X0_PGD N_A_c_363_n 5.17967e-19
cc_88 N_VDD_c_20_p N_A_c_363_n 4.32724e-19
cc_89 N_VDD_c_24_p N_A_c_363_n 4.10602e-19
cc_90 N_VDD_c_37_p N_A_c_363_n 4.1682e-19
cc_91 N_VDD_c_12_p N_A_c_363_n 3.91173e-19
cc_92 N_VDD_c_38_p N_A_c_363_n 5.53168e-19
cc_93 N_VDD_XI6.X0_S N_A_c_370_n 9.18655e-19
cc_94 N_VDD_c_12_p N_A_c_371_n 0.00608947f
cc_95 N_VDD_c_29_p N_A_c_372_n 8.16868e-19
cc_96 N_VDD_c_11_p N_A_c_372_n 2.36389e-19
cc_97 N_VDD_c_29_p N_A_c_374_n 6.33536e-19
cc_98 N_VDD_c_42_p N_A_c_374_n 5.39283e-19
cc_99 N_VDD_XI6.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_100 N_VDD_c_24_p N_BI_XI5.X0_D 3.7884e-19
cc_101 N_VDD_c_12_p N_BI_XI5.X0_D 3.48267e-19
cc_102 N_VDD_XI6.X0_S N_BI_c_443_n 3.48267e-19
cc_103 N_VDD_c_29_p N_BI_c_443_n 8.52765e-19
cc_104 N_VDD_c_24_p N_BI_c_443_n 4.58491e-19
cc_105 N_VDD_c_12_p N_BI_c_443_n 7.03408e-19
cc_106 N_VDD_c_24_p N_BI_c_447_n 2.4324e-19
cc_107 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_108 N_VDD_c_32_p N_AI_XI8.X0_D 3.73302e-19
cc_109 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.86706e-19
cc_110 N_VDD_c_110_p N_AI_c_513_n 2.86706e-19
cc_111 N_VDD_XI8.X0_S N_AI_c_514_n 3.48267e-19
cc_112 N_VDD_c_32_p N_AI_c_514_n 5.23123e-19
cc_113 N_VDD_c_20_p N_AI_c_514_n 5.01863e-19
cc_114 N_VDD_c_37_p N_AI_c_517_n 0.00111556f
cc_115 N_VDD_c_20_p N_AI_c_518_n 2.2965e-19
cc_116 N_VDD_XI9.X0_PGD N_B_XI5.X0_CG 9.5906e-19
cc_117 N_VDD_c_42_p N_B_XI5.X0_CG 9.74645e-19
cc_118 N_VDD_XI5.X0_PGD N_B_c_559_n 3.9688e-19
cc_119 N_VDD_XI7.X0_PGD N_B_c_559_n 2.07132e-19
cc_120 N_VDD_c_120_p N_B_c_561_n 9.5906e-19
cc_121 N_VDD_c_38_p N_B_c_562_n 2.92921e-19
cc_122 N_VDD_c_12_p N_B_c_563_n 5.34599e-19
cc_123 N_C_c_125_n N_VSS_XI10.X0_PGD 4.16623e-19
cc_124 N_C_c_136_p N_VSS_c_247_n 9.33417e-19
cc_125 C N_VSS_c_195_n 6.06998e-19
cc_126 N_C_c_138_p N_VSS_c_195_n 4.82229e-19
cc_127 N_C_c_139_p N_VSS_c_195_n 2.78014e-19
cc_128 N_C_c_138_p N_VSS_c_201_n 2.30642e-19
cc_129 N_C_c_133_n N_VSS_c_201_n 0.00197293f
cc_130 N_C_c_133_n N_VSS_c_209_n 0.00165406f
cc_131 N_C_c_143_p N_VSS_c_217_n 0.0041205f
cc_132 N_C_c_136_p N_VSS_c_217_n 7.00195e-19
cc_133 C N_VSS_c_217_n 4.56568e-19
cc_134 N_C_c_130_n N_VSS_c_217_n 6.1245e-19
cc_135 C N_VSS_c_228_n 2.17246e-19
cc_136 N_C_c_138_p N_VSS_c_228_n 4.01014e-19
cc_137 N_C_c_139_p N_VSS_c_228_n 4.34874e-19
cc_138 C N_VSS_c_233_n 2.70819e-19
cc_139 N_C_c_138_p N_VSS_c_233_n 9.65301e-19
cc_140 N_C_c_139_p N_VSS_c_233_n 0.00282977f
cc_141 N_C_c_133_n N_VSS_c_240_n 0.00175198f
cc_142 N_C_c_133_n N_CI_c_316_n 0.00136327f
cc_143 N_C_c_133_n N_CI_c_320_n 0.00242327f
cc_144 N_C_c_156_p N_CI_c_324_n 4.1018e-19
cc_145 N_C_c_133_n N_A_c_363_n 2.5075e-19
cc_146 N_C_c_158_p N_A_c_370_n 0.00148519f
cc_147 N_C_c_132_n N_A_c_370_n 8.20481e-19
cc_148 N_C_c_133_n N_A_c_370_n 2.96346e-19
cc_149 N_C_c_161_p N_A_c_370_n 2.4205e-19
cc_150 N_C_c_158_p N_A_c_381_n 0.00189731f
cc_151 N_C_c_132_n N_A_c_381_n 9.00742e-19
cc_152 N_C_c_133_n N_A_c_381_n 3.9734e-19
cc_153 N_C_c_156_p N_A_c_381_n 0.00207353f
cc_154 N_C_c_161_p N_A_c_381_n 6.32429e-19
cc_155 N_C_c_156_p N_A_c_386_n 5.4333e-19
cc_156 N_C_c_133_n N_BI_c_443_n 2.41407e-19
cc_157 N_C_c_133_n N_BI_c_447_n 4.13621e-19
cc_158 N_C_c_156_p N_BI_c_450_n 6.74177e-19
cc_159 N_C_c_156_p N_BI_c_451_n 0.00240592f
cc_160 N_C_c_158_p N_B_c_563_n 0.00168372f
cc_161 N_C_c_133_n N_B_c_563_n 0.0027048f
cc_162 N_C_c_156_p N_B_c_563_n 0.00182275f
cc_163 N_C_c_161_p N_B_c_563_n 2.1095e-19
cc_164 N_C_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_165 N_C_c_158_p N_Z_XI2.X0_D 3.48267e-19
cc_166 N_C_c_178_p N_Z_XI2.X0_D 3.48267e-19
cc_167 N_C_c_132_n N_Z_XI2.X0_D 3.43419e-19
cc_168 N_C_XI3.X0_S N_Z_c_624_n 3.48267e-19
cc_169 N_C_c_158_p N_Z_c_624_n 3.41702e-19
cc_170 N_C_c_178_p N_Z_c_624_n 5.7093e-19
cc_171 N_VSS_XI9.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_172 N_VSS_c_201_n N_CI_XI10.X0_D 3.48267e-19
cc_173 N_VSS_XI7.X0_S N_CI_XI4.X0_S 3.43419e-19
cc_174 N_VSS_c_213_n N_CI_XI4.X0_S 3.48267e-19
cc_175 N_VSS_XI9.X0_S N_CI_c_316_n 3.48267e-19
cc_176 N_VSS_c_195_n N_CI_c_316_n 5.78167e-19
cc_177 N_VSS_c_201_n N_CI_c_316_n 0.00107566f
cc_178 N_VSS_c_231_n N_CI_c_316_n 0.0020072f
cc_179 N_VSS_c_233_n N_CI_c_316_n 3.32126e-19
cc_180 N_VSS_XI7.X0_S N_CI_c_334_n 3.48267e-19
cc_181 N_VSS_c_213_n N_CI_c_334_n 9.13167e-19
cc_182 N_VSS_c_205_n N_CI_c_320_n 0.00134034f
cc_183 N_VSS_c_216_n N_CI_c_320_n 0.00393483f
cc_184 N_VSS_c_235_n N_CI_c_338_n 0.00292666f
cc_185 N_VSS_c_220_n N_A_c_387_n 0.00236445f
cc_186 N_VSS_XI8.X0_PGD N_A_c_362_n 3.86211e-19
cc_187 N_VSS_XI7.X0_S N_A_c_363_n 9.18655e-19
cc_188 N_VSS_c_213_n N_A_c_363_n 0.00149545f
cc_189 N_VSS_c_216_n N_A_c_363_n 2.12774e-19
cc_190 N_VSS_c_240_n N_A_c_363_n 2.27118e-19
cc_191 N_VSS_c_205_n N_A_c_372_n 4.58305e-19
cc_192 N_VSS_c_220_n N_A_c_372_n 4.30193e-19
cc_193 N_VSS_c_287_p N_A_c_374_n 8.53264e-19
cc_194 N_VSS_c_205_n N_A_c_374_n 4.26083e-19
cc_195 N_VSS_c_220_n N_A_c_374_n 7.20776e-19
cc_196 N_VSS_XI9.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_197 N_VSS_c_201_n N_BI_XI5.X0_D 3.48267e-19
cc_198 N_VSS_XI9.X0_S N_BI_c_443_n 3.48267e-19
cc_199 N_VSS_c_201_n N_BI_c_443_n 0.00102079f
cc_200 N_VSS_c_240_n N_BI_c_443_n 3.31365e-19
cc_201 N_VSS_c_216_n N_BI_c_457_n 2.90278e-19
cc_202 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_203 N_VSS_c_213_n N_AI_XI8.X0_D 3.48267e-19
cc_204 N_VSS_XI6.X0_PGD N_AI_XI2.X0_PGD 2.84687e-19
cc_205 N_VSS_c_213_n N_AI_XI2.X0_PGD 2.04949e-19
cc_206 N_VSS_c_192_n N_AI_c_523_n 2.84687e-19
cc_207 N_VSS_XI7.X0_S N_AI_c_514_n 3.48267e-19
cc_208 N_VSS_c_205_n N_AI_c_514_n 0.00163244f
cc_209 N_VSS_c_213_n N_AI_c_514_n 0.00129029f
cc_210 N_VSS_c_213_n N_AI_c_517_n 0.00168777f
cc_211 N_VSS_c_213_n N_AI_c_528_n 2.82216e-19
cc_212 N_VSS_c_216_n N_AI_c_518_n 0.00857137f
cc_213 N_VSS_c_224_n N_B_XI6.X0_CG 0.00272012f
cc_214 N_VSS_XI8.X0_PGD N_B_c_559_n 2.07132e-19
cc_215 N_VSS_XI6.X0_PGD N_B_c_559_n 3.923e-19
cc_216 N_VSS_c_224_n N_B_c_571_n 0.00138168f
cc_217 N_VSS_c_209_n B 5.92764e-19
cc_218 N_VSS_c_224_n N_B_c_562_n 6.1245e-19
cc_219 N_VSS_c_209_n N_B_c_563_n 6.44904e-19
cc_220 N_CI_c_316_n N_BI_c_443_n 0.00104494f
cc_221 N_CI_c_324_n N_BI_c_459_n 6.86101e-19
cc_222 N_CI_c_334_n N_BI_c_447_n 8.7e-19
cc_223 N_CI_c_320_n N_BI_c_447_n 9.27611e-19
cc_224 N_CI_c_324_n N_BI_c_450_n 0.00228179f
cc_225 N_CI_c_316_n N_AI_c_514_n 5.24832e-19
cc_226 N_CI_c_334_n N_AI_c_514_n 5.10362e-19
cc_227 N_CI_c_334_n N_AI_c_517_n 0.00202744f
cc_228 N_CI_c_320_n N_AI_c_517_n 0.00654866f
cc_229 N_CI_c_324_n N_AI_c_517_n 0.00288502f
cc_230 N_CI_c_349_p N_AI_c_517_n 8.49574e-19
cc_231 N_CI_c_320_n N_AI_c_518_n 9.37419e-19
cc_232 N_CI_c_324_n N_B_c_575_n 0.00103435f
cc_233 N_CI_c_324_n N_B_c_576_n 2.42418e-19
cc_234 N_CI_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_235 N_CI_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_236 N_CI_c_334_n N_Z_XI4.X0_D 3.48267e-19
cc_237 N_CI_c_356_p N_Z_XI4.X0_D 3.48267e-19
cc_238 N_CI_XI4.X0_S N_Z_c_624_n 3.48267e-19
cc_239 N_CI_XI1.X0_S N_Z_c_624_n 3.48267e-19
cc_240 N_CI_c_334_n N_Z_c_624_n 5.68744e-19
cc_241 N_CI_c_356_p N_Z_c_624_n 5.68744e-19
cc_242 N_A_XI3.X0_PGD N_BI_XI3.X0_CG 8.79767e-19
cc_243 N_A_c_399_p N_BI_XI3.X0_CG 0.00237738f
cc_244 N_A_c_399_p N_BI_c_465_n 0.00117691f
cc_245 N_A_c_363_n N_BI_c_443_n 4.0484e-19
cc_246 N_A_c_370_n N_BI_c_443_n 6.63236e-19
cc_247 N_A_c_363_n N_BI_c_468_n 2.37396e-19
cc_248 N_A_c_386_n N_BI_c_459_n 7.92141e-19
cc_249 N_A_c_399_p N_BI_c_459_n 4.87897e-19
cc_250 N_A_c_363_n N_BI_c_471_n 3.8563e-19
cc_251 N_A_XI3.X0_PGD N_BI_c_472_n 0.00133285f
cc_252 N_A_c_386_n N_BI_c_472_n 4.79282e-19
cc_253 N_A_c_399_p N_BI_c_472_n 0.00152548f
cc_254 N_A_c_370_n N_BI_c_447_n 0.00181644f
cc_255 N_A_c_363_n N_BI_c_457_n 0.00247154f
cc_256 N_A_c_370_n N_BI_c_477_n 2.27623e-19
cc_257 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174824f
cc_258 N_A_c_370_n N_AI_XI2.X0_PGD 8.597e-19
cc_259 N_A_c_415_p N_AI_c_523_n 0.00199346f
cc_260 N_A_c_381_n N_AI_c_523_n 0.00123218f
cc_261 N_A_c_417_p N_AI_c_513_n 0.00202303f
cc_262 N_A_c_363_n N_AI_c_514_n 0.00165136f
cc_263 N_A_c_363_n N_AI_c_517_n 0.00184834f
cc_264 N_A_c_362_n N_B_c_559_n 0.00360254f
cc_265 N_A_c_363_n N_B_c_559_n 5.41329e-19
cc_266 N_A_c_374_n N_B_c_561_n 4.14098e-19
cc_267 N_A_c_381_n N_B_c_580_n 2.74862e-19
cc_268 N_A_XI3.X0_PGD N_B_c_581_n 8.79767e-19
cc_269 N_A_c_363_n B 6.972e-19
cc_270 N_A_c_370_n B 3.89684e-19
cc_271 N_A_c_370_n N_B_c_584_n 3.55503e-19
cc_272 N_A_c_381_n N_B_c_584_n 4.94081e-19
cc_273 N_A_c_381_n N_B_c_575_n 3.26384e-19
cc_274 N_A_c_362_n N_B_c_562_n 2.86506e-19
cc_275 N_A_c_370_n N_B_c_562_n 6.34732e-19
cc_276 N_A_c_370_n N_B_c_589_n 3.37713e-19
cc_277 N_A_XI3.X0_PGD N_B_c_590_n 0.00133285f
cc_278 N_A_c_370_n N_B_c_563_n 0.00206097f
cc_279 N_A_c_381_n N_B_c_563_n 0.00238641f
cc_280 N_A_c_381_n N_Z_XI2.X0_D 6.94686e-19
cc_281 N_A_XI3.X0_PGD N_Z_c_624_n 6.45939e-19
cc_282 N_A_c_370_n N_Z_c_624_n 0.00131646f
cc_283 N_A_c_381_n N_Z_c_624_n 0.00121415f
cc_284 N_BI_c_478_p N_AI_XI2.X0_PGD 8.79767e-19
cc_285 N_BI_c_471_n N_AI_XI2.X0_PGD 0.00133285f
cc_286 N_BI_c_471_n N_AI_c_546_n 6.37981e-19
cc_287 N_BI_c_457_n N_AI_c_514_n 8.05284e-19
cc_288 N_BI_c_468_n N_AI_c_517_n 4.93364e-19
cc_289 N_BI_c_447_n N_AI_c_517_n 0.00402897f
cc_290 N_BI_c_477_n N_AI_c_517_n 4.42808e-19
cc_291 N_BI_c_478_p N_AI_c_528_n 0.00234569f
cc_292 N_BI_c_468_n N_AI_c_528_n 4.6759e-19
cc_293 N_BI_c_471_n N_AI_c_528_n 0.00166302f
cc_294 N_BI_c_443_n B 4.30856e-19
cc_295 N_BI_c_447_n B 3.14738e-19
cc_296 N_BI_c_468_n N_B_c_584_n 5.92939e-19
cc_297 N_BI_c_477_n N_B_c_584_n 3.24098e-19
cc_298 N_BI_c_459_n N_B_c_575_n 0.0018551f
cc_299 N_BI_c_471_n N_B_c_589_n 0.00266367f
cc_300 N_BI_c_472_n N_B_c_589_n 6.17967e-19
cc_301 N_BI_c_471_n N_B_c_590_n 7.16621e-19
cc_302 N_BI_c_472_n N_B_c_590_n 0.00243799f
cc_303 N_BI_c_443_n N_B_c_563_n 0.00165434f
cc_304 N_BI_c_459_n N_B_c_563_n 0.00159414f
cc_305 N_BI_c_447_n N_B_c_563_n 0.0157983f
cc_306 N_BI_c_450_n N_B_c_563_n 6.88876e-19
cc_307 N_BI_c_451_n N_B_c_563_n 8.27361e-19
cc_308 N_BI_c_477_n N_B_c_607_n 0.00346365f
cc_309 N_BI_c_503_p N_B_c_607_n 0.00194674f
cc_310 N_BI_c_468_n N_B_c_576_n 3.02576e-19
cc_311 N_BI_c_450_n N_B_c_576_n 8.19447e-19
cc_312 N_BI_c_468_n N_Z_c_624_n 0.00155391f
cc_313 N_BI_c_459_n N_Z_c_624_n 0.00136914f
cc_314 N_BI_c_472_n N_Z_c_624_n 8.66889e-19
cc_315 N_BI_c_477_n N_Z_c_624_n 4.81308e-19
cc_316 N_AI_XI2.X0_PGD N_B_XI2.X0_CG 8.63152e-19
cc_317 N_AI_XI2.X0_PGD N_B_c_589_n 0.00133285f
cc_318 N_AI_XI2.X0_PGD N_Z_c_624_n 3.30612e-19
cc_319 N_B_c_584_n N_Z_c_624_n 0.00130267f
cc_320 N_B_c_575_n N_Z_c_624_n 0.00130267f
cc_321 N_B_c_589_n N_Z_c_624_n 8.66889e-19
cc_322 N_B_c_590_n N_Z_c_624_n 8.66889e-19
cc_323 N_B_c_563_n N_Z_c_624_n 0.00103251f
cc_324 N_B_c_607_n N_Z_c_624_n 0.00216955f
cc_325 N_B_c_576_n N_Z_c_624_n 9.92382e-19
*
.ends
*
*
.subckt XNOR3_HPNW4 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XNOR3_N1_2
.ends
*
* File: G4_XOR2_N1.pex.netlist
* Created: Fri Mar 18 15:34:38 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*







.subckt G4_XOR2_N1_2 VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI1.X0 N_NET1_XI1.X0_D N_VDD_XI1.X0_PGD N_B_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI9.X0 N_NET2_XI9.X0_D N_VSS_XI9.X0_PGD N_A_XI9.X0_CG N_VSS_XI9.X0_PGD
+ N_VDD_XI9.X0_S TIGFET_HPNW4
XI10.X0 N_NET1_XI1.X0_D N_VSS_XI10.X0_PGD N_B_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW4
XI3.X0 N_NET2_XI9.X0_D N_VDD_XI3.X0_PGD N_A_XI3.X0_CG N_VDD_XI3.X0_PGD
+ N_VSS_XI3.X0_S TIGFET_HPNW4
XI5.X0 N_Z_XI5.X0_D N_B_XI5.X0_PGD N_NET2_XI5.X0_CG N_B_XI5.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW4
XI8.X0 N_Z_XI8.X0_D N_A_XI8.X0_PGD N_B_XI8.X0_CG N_A_XI8.X0_PGD N_VSS_XI3.X0_S
+ TIGFET_HPNW4
XI11.X0 N_Z_XI5.X0_D N_NET1_XI11.X0_PGD N_A_XI11.X0_CG N_NET1_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW4
XI7.X0 N_Z_XI8.X0_D N_NET2_XI7.X0_PGD N_NET1_XI7.X0_CG N_NET2_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW4
*
x_PM_G4_XOR2_N1_VSS N_VSS_XI1.X0_S N_VSS_XI9.X0_PGD N_VSS_XI10.X0_PGD
+ N_VSS_XI3.X0_S N_VSS_XI7.X0_S N_VSS_c_8_p N_VSS_c_23_p N_VSS_c_56_p
+ N_VSS_c_40_p N_VSS_c_7_p N_VSS_c_3_p N_VSS_c_13_p N_VSS_c_30_p N_VSS_c_4_p
+ N_VSS_c_6_p N_VSS_c_14_p N_VSS_c_31_p N_VSS_c_10_p N_VSS_c_11_p N_VSS_c_18_p
+ N_VSS_c_19_p N_VSS_c_26_p N_VSS_c_29_p N_VSS_c_27_p N_VSS_c_62_p N_VSS_c_46_p
+ N_VSS_c_83_p N_VSS_c_12_p N_VSS_c_28_p VSS Vss PM_G4_XOR2_N1_VSS
x_PM_G4_XOR2_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI9.X0_S N_VDD_XI10.X0_S
+ N_VDD_XI3.X0_PGD N_VDD_XI11.X0_S N_VDD_c_112_n N_VDD_c_163_p N_VDD_c_113_n
+ N_VDD_c_114_n N_VDD_c_118_n N_VDD_c_121_n N_VDD_c_124_n N_VDD_c_125_n
+ N_VDD_c_127_n N_VDD_c_134_n N_VDD_c_135_n N_VDD_c_137_n N_VDD_c_141_n
+ N_VDD_c_144_n N_VDD_c_168_p N_VDD_c_149_n N_VDD_c_182_p N_VDD_c_152_n
+ N_VDD_c_153_n VDD N_VDD_c_154_n N_VDD_c_156_n Vss PM_G4_XOR2_N1_VDD
x_PM_G4_XOR2_N1_A N_A_XI9.X0_CG N_A_XI3.X0_CG N_A_XI8.X0_PGD N_A_XI11.X0_CG
+ N_A_c_212_n N_A_c_213_n N_A_c_215_n N_A_c_216_n N_A_c_246_p N_A_c_231_n A
+ N_A_c_219_n N_A_c_223_n N_A_c_224_n N_A_c_239_n N_A_c_242_p N_A_c_240_n Vss
+ PM_G4_XOR2_N1_A
x_PM_G4_XOR2_N1_NET1 N_NET1_XI1.X0_D N_NET1_XI11.X0_PGD N_NET1_XI7.X0_CG
+ N_NET1_c_282_n N_NET1_c_302_p N_NET1_c_273_n N_NET1_c_276_n N_NET1_c_289_n
+ N_NET1_c_277_n Vss PM_G4_XOR2_N1_NET1
x_PM_G4_XOR2_N1_NET2 N_NET2_XI9.X0_D N_NET2_XI5.X0_CG N_NET2_XI7.X0_PGD
+ N_NET2_c_333_n N_NET2_c_352_p N_NET2_c_334_n N_NET2_c_335_n N_NET2_c_314_n
+ N_NET2_c_318_n N_NET2_c_338_n N_NET2_c_321_n Vss PM_G4_XOR2_N1_NET2
x_PM_G4_XOR2_N1_B N_B_XI1.X0_CG N_B_XI10.X0_CG N_B_XI5.X0_PGD N_B_XI8.X0_CG
+ N_B_c_360_n N_B_c_381_n N_B_c_362_n N_B_c_363_n N_B_c_392_n N_B_c_364_n
+ N_B_c_393_n N_B_c_383_n B N_B_c_365_n N_B_c_367_n Vss PM_G4_XOR2_N1_B
x_PM_G4_XOR2_N1_Z N_Z_XI5.X0_D N_Z_XI8.X0_D N_Z_c_401_n Z Vss PM_G4_XOR2_N1_Z
cc_1 N_VSS_XI9.X0_PGD N_VDD_XI1.X0_PGD 2.77144e-19
cc_2 N_VSS_XI10.X0_PGD N_VDD_XI1.X0_PGD 0.00167677f
cc_3 N_VSS_c_3_p N_VDD_XI9.X0_S 2.05974e-19
cc_4 N_VSS_c_4_p N_VDD_XI10.X0_S 2.02468e-19
cc_5 N_VSS_XI9.X0_PGD N_VDD_XI3.X0_PGD 0.00169392f
cc_6 N_VSS_c_6_p N_VDD_XI11.X0_S 2.02468e-19
cc_7 N_VSS_c_7_p N_VDD_c_112_n 0.00167677f
cc_8 N_VSS_c_8_p N_VDD_c_113_n 0.00169392f
cc_9 N_VSS_c_3_p N_VDD_c_114_n 0.00187494f
cc_10 N_VSS_c_10_p N_VDD_c_114_n 0.00305883f
cc_11 N_VSS_c_11_p N_VDD_c_114_n 0.00593001f
cc_12 N_VSS_c_12_p N_VDD_c_114_n 8.91588e-19
cc_13 N_VSS_c_13_p N_VDD_c_118_n 4.43871e-19
cc_14 N_VSS_c_14_p N_VDD_c_118_n 3.66936e-19
cc_15 N_VSS_c_11_p N_VDD_c_118_n 0.0030181f
cc_16 N_VSS_XI1.X0_S N_VDD_c_121_n 3.7884e-19
cc_17 N_VSS_c_3_p N_VDD_c_121_n 4.73473e-19
cc_18 N_VSS_c_18_p N_VDD_c_121_n 0.00352628f
cc_19 N_VSS_c_19_p N_VDD_c_124_n 0.0010586f
cc_20 N_VSS_XI1.X0_S N_VDD_c_125_n 2.02468e-19
cc_21 N_VSS_c_3_p N_VDD_c_125_n 8.57018e-19
cc_22 N_VSS_c_8_p N_VDD_c_127_n 3.60588e-19
cc_23 N_VSS_c_23_p N_VDD_c_127_n 3.60588e-19
cc_24 N_VSS_c_13_p N_VDD_c_127_n 0.00141228f
cc_25 N_VSS_c_14_p N_VDD_c_127_n 0.00112249f
cc_26 N_VSS_c_26_p N_VDD_c_127_n 0.00343125f
cc_27 N_VSS_c_27_p N_VDD_c_127_n 0.0059942f
cc_28 N_VSS_c_28_p N_VDD_c_127_n 7.74609e-19
cc_29 N_VSS_c_29_p N_VDD_c_134_n 0.00107456f
cc_30 N_VSS_c_30_p N_VDD_c_135_n 9.22488e-19
cc_31 N_VSS_c_31_p N_VDD_c_135_n 3.82294e-19
cc_32 N_VSS_c_7_p N_VDD_c_137_n 3.60588e-19
cc_33 N_VSS_c_30_p N_VDD_c_137_n 0.00161703f
cc_34 N_VSS_c_31_p N_VDD_c_137_n 2.03837e-19
cc_35 N_VSS_c_18_p N_VDD_c_137_n 0.00605426f
cc_36 N_VSS_c_13_p N_VDD_c_141_n 9.25616e-19
cc_37 N_VSS_c_4_p N_VDD_c_141_n 9.18823e-19
cc_38 N_VSS_c_14_p N_VDD_c_141_n 3.99794e-19
cc_39 N_VSS_XI3.X0_S N_VDD_c_144_n 2.21516e-19
cc_40 N_VSS_c_40_p N_VDD_c_144_n 2.69489e-19
cc_41 N_VSS_c_30_p N_VDD_c_144_n 0.0023129f
cc_42 N_VSS_c_4_p N_VDD_c_144_n 2.43341e-19
cc_43 N_VSS_c_31_p N_VDD_c_144_n 9.55109e-19
cc_44 N_VSS_XI7.X0_S N_VDD_c_149_n 2.02468e-19
cc_45 N_VSS_c_6_p N_VDD_c_149_n 2.98086e-19
cc_46 N_VSS_c_46_p N_VDD_c_149_n 0.00130737f
cc_47 N_VSS_c_11_p N_VDD_c_152_n 9.23211e-19
cc_48 N_VSS_c_18_p N_VDD_c_153_n 0.0010761f
cc_49 N_VSS_c_30_p N_VDD_c_154_n 3.48267e-19
cc_50 N_VSS_c_31_p N_VDD_c_154_n 8.0279e-19
cc_51 N_VSS_c_13_p N_VDD_c_156_n 3.48267e-19
cc_52 N_VSS_c_14_p N_VDD_c_156_n 8.07896e-19
cc_53 N_VSS_c_14_p N_A_c_212_n 0.00234108f
cc_54 N_VSS_XI9.X0_PGD N_A_c_213_n 3.99472e-19
cc_55 N_VSS_XI10.X0_PGD N_A_c_213_n 2.20169e-19
cc_56 N_VSS_c_56_p N_A_c_215_n 9.41527e-19
cc_57 N_VSS_XI10.X0_PGD N_A_c_216_n 2.20169e-19
cc_58 N_VSS_c_13_p A 5.59945e-19
cc_59 N_VSS_c_14_p A 4.56568e-19
cc_60 N_VSS_c_4_p N_A_c_219_n 0.00506909f
cc_61 N_VSS_c_11_p N_A_c_219_n 6.18143e-19
cc_62 N_VSS_c_62_p N_A_c_219_n 0.00198136f
cc_63 N_VSS_c_46_p N_A_c_219_n 2.97351e-19
cc_64 N_VSS_c_62_p N_A_c_223_n 0.00118029f
cc_65 N_VSS_c_13_p N_A_c_224_n 4.56568e-19
cc_66 N_VSS_c_14_p N_A_c_224_n 6.1245e-19
cc_67 N_VSS_XI1.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_68 N_VSS_c_3_p N_NET1_XI1.X0_D 3.48267e-19
cc_69 N_VSS_XI1.X0_S N_NET1_c_273_n 3.48267e-19
cc_70 N_VSS_c_3_p N_NET1_c_273_n 0.00108327f
cc_71 N_VSS_c_18_p N_NET1_c_273_n 3.32126e-19
cc_72 N_VSS_c_30_p N_NET1_c_276_n 0.00167316f
cc_73 N_VSS_c_10_p N_NET1_c_277_n 3.27829e-19
cc_74 N_VSS_c_18_p N_NET1_c_277_n 6.3226e-19
cc_75 N_VSS_XI3.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_76 N_VSS_c_4_p N_NET2_XI9.X0_D 3.48267e-19
cc_77 N_VSS_XI3.X0_S N_NET2_c_314_n 3.48267e-19
cc_78 N_VSS_c_4_p N_NET2_c_314_n 0.00151106f
cc_79 N_VSS_c_11_p N_NET2_c_314_n 5.08641e-19
cc_80 N_VSS_c_27_p N_NET2_c_314_n 3.31434e-19
cc_81 N_VSS_c_4_p N_NET2_c_318_n 0.00228146f
cc_82 N_VSS_c_62_p N_NET2_c_318_n 0.00565735f
cc_83 N_VSS_c_83_p N_NET2_c_318_n 0.00115259f
cc_84 N_VSS_c_13_p N_NET2_c_321_n 5.79036e-19
cc_85 N_VSS_c_27_p N_NET2_c_321_n 0.00176418f
cc_86 N_VSS_c_31_p N_B_XI10.X0_CG 0.00234108f
cc_87 N_VSS_XI10.X0_PGD N_B_XI5.X0_PGD 0.00176522f
cc_88 N_VSS_XI9.X0_PGD N_B_c_360_n 2.20169e-19
cc_89 N_VSS_XI10.X0_PGD N_B_c_360_n 3.99472e-19
cc_90 N_VSS_XI10.X0_PGD N_B_c_362_n 4.05198e-19
cc_91 N_VSS_c_31_p N_B_c_363_n 9.49637e-19
cc_92 N_VSS_c_40_p N_B_c_364_n 0.00154836f
cc_93 N_VSS_c_30_p N_B_c_365_n 5.01474e-19
cc_94 N_VSS_c_31_p N_B_c_365_n 4.56568e-19
cc_95 N_VSS_c_30_p N_B_c_367_n 4.56568e-19
cc_96 N_VSS_c_31_p N_B_c_367_n 6.1245e-19
cc_97 N_VSS_XI3.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_98 N_VSS_XI7.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_99 N_VSS_c_4_p N_Z_XI8.X0_D 3.48267e-19
cc_100 N_VSS_c_6_p N_Z_XI8.X0_D 3.48267e-19
cc_101 N_VSS_XI3.X0_S N_Z_c_401_n 3.48267e-19
cc_102 N_VSS_XI7.X0_S N_Z_c_401_n 3.48267e-19
cc_103 N_VSS_c_4_p N_Z_c_401_n 4.94062e-19
cc_104 N_VSS_c_6_p N_Z_c_401_n 5.68744e-19
cc_105 N_VSS_c_62_p N_Z_c_401_n 3.25705e-19
cc_106 N_VDD_c_156_n N_A_XI3.X0_CG 9.28877e-19
cc_107 N_VDD_XI3.X0_PGD N_A_XI8.X0_PGD 0.00157721f
cc_108 N_VDD_XI1.X0_PGD N_A_c_213_n 2.20169e-19
cc_109 N_VDD_XI3.X0_PGD N_A_c_213_n 4.04053e-19
cc_110 N_VDD_XI3.X0_PGD N_A_c_216_n 4.05198e-19
cc_111 N_VDD_c_163_p N_A_c_231_n 0.00157721f
cc_112 N_VDD_c_114_n A 3.46645e-19
cc_113 N_VDD_c_135_n A 2.52205e-19
cc_114 N_VDD_c_141_n N_A_c_219_n 5.08705e-19
cc_115 N_VDD_c_156_n N_A_c_219_n 3.5189e-19
cc_116 N_VDD_c_168_p N_A_c_223_n 8.44396e-19
cc_117 N_VDD_c_114_n N_A_c_224_n 4.71537e-19
cc_118 N_VDD_c_154_n N_A_c_224_n 4.4222e-19
cc_119 N_VDD_c_156_n N_A_c_239_n 9.06702e-19
cc_120 N_VDD_c_168_p N_A_c_240_n 0.00102412f
cc_121 N_VDD_XI10.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_122 N_VDD_c_137_n N_NET1_XI1.X0_D 3.7884e-19
cc_123 N_VDD_c_144_n N_NET1_XI1.X0_D 3.48267e-19
cc_124 N_VDD_c_168_p N_NET1_c_282_n 8.23105e-19
cc_125 N_VDD_XI10.X0_S N_NET1_c_273_n 3.48267e-19
cc_126 N_VDD_c_137_n N_NET1_c_273_n 4.58491e-19
cc_127 N_VDD_c_144_n N_NET1_c_273_n 0.00110118f
cc_128 N_VDD_c_144_n N_NET1_c_276_n 0.00124814f
cc_129 N_VDD_c_168_p N_NET1_c_276_n 0.00341061f
cc_130 N_VDD_c_182_p N_NET1_c_276_n 8.21148e-19
cc_131 N_VDD_c_144_n N_NET1_c_289_n 2.78343e-19
cc_132 N_VDD_c_168_p N_NET1_c_289_n 0.00115624f
cc_133 N_VDD_c_182_p N_NET1_c_289_n 3.70842e-19
cc_134 N_VDD_c_135_n N_NET1_c_277_n 2.90608e-19
cc_135 N_VDD_XI9.X0_S N_NET2_XI9.X0_D 3.67949e-19
cc_136 N_VDD_c_125_n N_NET2_XI9.X0_D 3.72199e-19
cc_137 N_VDD_XI9.X0_S N_NET2_c_314_n 3.9802e-19
cc_138 N_VDD_c_125_n N_NET2_c_314_n 5.226e-19
cc_139 N_VDD_c_127_n N_NET2_c_314_n 5.01863e-19
cc_140 N_VDD_c_141_n N_NET2_c_318_n 2.9893e-19
cc_141 N_VDD_c_114_n N_B_XI1.X0_CG 3.37985e-19
cc_142 N_VDD_c_154_n N_B_XI1.X0_CG 9.28877e-19
cc_143 N_VDD_XI1.X0_PGD N_B_c_360_n 4.04053e-19
cc_144 N_VDD_XI3.X0_PGD N_B_c_360_n 2.20169e-19
cc_145 N_VDD_XI3.X0_PGD N_B_c_362_n 2.20169e-19
cc_146 N_VDD_c_144_n N_B_c_364_n 2.75901e-19
cc_147 N_VDD_c_168_p N_B_c_364_n 9.79508e-19
cc_148 N_VDD_c_141_n N_B_c_365_n 2.10322e-19
cc_149 N_VDD_c_156_n N_B_c_367_n 4.24849e-19
cc_150 N_VDD_XI10.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_151 N_VDD_XI11.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_152 N_VDD_c_144_n N_Z_XI5.X0_D 3.48267e-19
cc_153 N_VDD_c_168_p N_Z_XI5.X0_D 3.7884e-19
cc_154 N_VDD_c_149_n N_Z_XI5.X0_D 3.72199e-19
cc_155 N_VDD_XI10.X0_S N_Z_c_401_n 3.48267e-19
cc_156 N_VDD_XI11.X0_S N_Z_c_401_n 3.48267e-19
cc_157 N_VDD_c_144_n N_Z_c_401_n 7.90262e-19
cc_158 N_VDD_c_168_p N_Z_c_401_n 6.5261e-19
cc_159 N_VDD_c_149_n N_Z_c_401_n 8.53368e-19
cc_160 N_A_XI11.X0_CG N_NET1_XI11.X0_PGD 4.5346e-19
cc_161 N_A_c_242_p N_NET1_XI11.X0_PGD 0.0013363f
cc_162 N_A_c_223_n N_NET1_c_276_n 0.00121138f
cc_163 N_A_c_240_n N_NET1_c_276_n 0.00197573f
cc_164 N_A_XI11.X0_CG N_NET1_c_289_n 0.00234108f
cc_165 N_A_c_246_p N_NET1_c_289_n 0.00110158f
cc_166 N_A_c_242_p N_NET1_c_289_n 0.0014909f
cc_167 N_A_c_242_p N_NET2_XI5.X0_CG 2.18475e-19
cc_168 N_A_XI8.X0_PGD N_NET2_XI7.X0_PGD 0.00161543f
cc_169 N_A_c_216_n N_NET2_XI7.X0_PGD 3.14428e-19
cc_170 N_A_c_242_p N_NET2_XI7.X0_PGD 4.01857e-19
cc_171 N_A_XI8.X0_PGD N_NET2_c_333_n 4.60549e-19
cc_172 N_A_c_246_p N_NET2_c_334_n 2.17364e-19
cc_173 N_A_c_231_n N_NET2_c_335_n 0.00161543f
cc_174 N_A_c_219_n N_NET2_c_318_n 0.00221613f
cc_175 N_A_c_223_n N_NET2_c_318_n 7.30894e-19
cc_176 N_A_c_219_n N_NET2_c_338_n 3.44698e-19
cc_177 N_A_c_239_n N_NET2_c_338_n 9.17176e-19
cc_178 N_A_c_242_p N_NET2_c_338_n 3.34137e-19
cc_179 N_A_c_216_n N_B_XI8.X0_CG 0.003858f
cc_180 N_A_c_239_n N_B_XI8.X0_CG 0.00111269f
cc_181 N_A_c_213_n N_B_c_360_n 0.00504555f
cc_182 N_A_c_224_n N_B_c_381_n 3.67702e-19
cc_183 N_A_c_216_n N_B_c_362_n 0.00373351f
cc_184 N_A_c_216_n N_B_c_383_n 0.00215664f
cc_185 N_A_c_240_n N_B_c_365_n 2.66007e-19
cc_186 N_A_c_213_n N_B_c_367_n 4.25664e-19
cc_187 N_A_c_219_n N_Z_c_401_n 0.00323423f
cc_188 N_A_c_223_n N_Z_c_401_n 0.00319047f
cc_189 N_A_c_242_p N_Z_c_401_n 8.50872e-19
cc_190 N_NET1_c_273_n N_NET2_XI9.X0_D 2.02468e-19
cc_191 N_NET1_XI11.X0_PGD N_NET2_XI5.X0_CG 3.25363e-19
cc_192 N_NET1_c_302_p N_NET2_XI7.X0_PGD 0.00868439f
cc_193 N_NET1_XI11.X0_PGD N_NET2_c_333_n 0.00320236f
cc_194 N_NET1_XI1.X0_D N_NET2_c_314_n 2.02468e-19
cc_195 N_NET1_c_273_n N_NET2_c_314_n 3.48409e-19
cc_196 N_NET1_c_276_n N_NET2_c_318_n 0.00270459f
cc_197 N_NET1_XI7.X0_CG N_NET2_c_338_n 0.00266268f
cc_198 N_NET1_XI11.X0_PGD N_B_XI5.X0_PGD 0.00188194f
cc_199 N_NET1_XI7.X0_CG N_B_XI8.X0_CG 2.72153e-19
cc_200 N_NET1_c_282_n N_B_c_364_n 0.00165596f
cc_201 N_NET1_c_302_p N_B_c_383_n 2.72153e-19
cc_202 N_NET2_XI5.X0_CG N_B_XI5.X0_PGD 0.00233046f
cc_203 N_NET2_c_333_n N_B_XI5.X0_PGD 0.00159876f
cc_204 N_NET2_XI7.X0_PGD N_B_c_392_n 4.0517e-19
cc_205 N_NET2_c_352_p N_B_c_393_n 0.00233046f
cc_206 N_NET2_XI7.X0_PGD N_B_c_383_n 0.00313315f
cc_207 N_NET2_c_352_p N_B_c_383_n 0.00171842f
cc_208 N_NET2_XI7.X0_PGD N_Z_c_401_n 0.0012119f
cc_209 N_NET2_c_333_n N_Z_c_401_n 4.14549e-19
cc_210 N_NET2_c_318_n N_Z_c_401_n 2.62894e-19
cc_211 N_B_c_383_n N_Z_c_401_n 8.74847e-19
*
.ends
*
*
.subckt XOR2_HPNW4 A B Y VDD VSS
xgate (VSS VDD A B Y) G4_XOR2_N1_2
.ends
*
* File: G5_XOR3_N1.pex.netlist
* Created: Sun Apr 10 19:25:53 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*









.subckt G5_XOR3_N1_2 VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI10.X0 N_CI_XI10.X0_D N_VSS_XI10.X0_PGD N_C_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW4
XI9.X0 N_CI_XI10.X0_D N_VDD_XI9.X0_PGD N_C_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI5.X0 N_BI_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI6.X0 N_BI_XI5.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW4
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW4
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_BI_XI2.X0_CG N_AI_XI2.X0_PGD N_C_XI2.X0_S
+ TIGFET_HPNW4
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_B_XI4.X0_CG N_AI_XI4.X0_PGD N_CI_XI4.X0_S
+ TIGFET_HPNW4
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_B_XI3.X0_CG N_A_XI3.X0_PGD N_C_XI3.X0_S
+ TIGFET_HPNW4
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_BI_XI1.X0_CG N_A_XI1.X0_PGD N_CI_XI1.X0_S
+ TIGFET_HPNW4
*
x_PM_G5_XOR3_N1_VDD N_VDD_XI10.X0_S N_VDD_XI9.X0_PGD N_VDD_XI5.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI6.X0_S N_VDD_XI7.X0_PGD N_VDD_c_121_p N_VDD_c_20_p
+ N_VDD_c_25_p N_VDD_c_4_p N_VDD_c_109_p N_VDD_c_21_p N_VDD_c_6_p N_VDD_c_27_p
+ N_VDD_c_5_p N_VDD_c_64_p N_VDD_c_29_p N_VDD_c_30_p N_VDD_c_31_p N_VDD_c_37_p
+ N_VDD_c_34_p N_VDD_c_22_p N_VDD_c_11_p N_VDD_c_26_p N_VDD_c_39_p N_VDD_c_12_p
+ N_VDD_c_60_p VDD N_VDD_c_68_p N_VDD_c_72_p N_VDD_c_19_p N_VDD_c_2_p
+ N_VDD_c_44_p N_VDD_c_40_p Vss PM_G5_XOR3_N1_VDD
x_PM_G5_XOR3_N1_C N_C_XI10.X0_CG N_C_XI9.X0_CG N_C_XI2.X0_S N_C_XI3.X0_S
+ N_C_c_144_p N_C_c_127_n C N_C_c_140_p N_C_c_157_p N_C_c_179_p N_C_c_132_n
+ N_C_c_134_n N_C_c_135_n N_C_c_156_p N_C_c_141_p N_C_c_160_p Vss
+ PM_G5_XOR3_N1_C
x_PM_G5_XOR3_N1_VSS N_VSS_XI10.X0_PGD N_VSS_XI9.X0_S N_VSS_XI8.X0_PGD
+ N_VSS_XI6.X0_PGD N_VSS_XI7.X0_S N_VSS_c_191_n N_VSS_c_250_n N_VSS_c_192_n
+ N_VSS_c_194_n N_VSS_c_288_p N_VSS_c_195_n N_VSS_c_196_n N_VSS_c_198_n
+ N_VSS_c_204_n N_VSS_c_208_n N_VSS_c_212_n N_VSS_c_216_n N_VSS_c_218_n
+ N_VSS_c_221_n N_VSS_c_225_n N_VSS_c_229_n N_VSS_c_232_n N_VSS_c_234_n
+ N_VSS_c_235_n N_VSS_c_236_n N_VSS_c_240_n N_VSS_c_241_n N_VSS_c_244_n VSS
+ N_VSS_c_246_n N_VSS_c_247_n N_VSS_c_248_n Vss PM_G5_XOR3_N1_VSS
x_PM_G5_XOR3_N1_CI N_CI_XI10.X0_D N_CI_XI4.X0_S N_CI_XI1.X0_S N_CI_c_317_n
+ N_CI_c_333_n N_CI_c_373_p N_CI_c_321_n N_CI_c_337_n N_CI_c_339_n N_CI_c_347_p
+ N_CI_c_356_p N_CI_c_325_n Vss PM_G5_XOR3_N1_CI
x_PM_G5_XOR3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI3.X0_PGD N_A_XI1.X0_PGD
+ N_A_c_402_n N_A_c_378_n N_A_c_428_p N_A_c_430_p N_A_c_379_n N_A_c_387_n
+ N_A_c_396_n N_A_c_388_n A N_A_c_389_n N_A_c_401_n N_A_c_390_n N_A_c_434_p Vss
+ PM_G5_XOR3_N1_A
x_PM_G5_XOR3_N1_BI N_BI_XI5.X0_D N_BI_XI2.X0_CG N_BI_XI1.X0_CG N_BI_c_480_n
+ N_BI_c_481_n N_BI_c_460_n N_BI_c_464_n N_BI_c_478_n N_BI_c_486_n N_BI_c_487_n
+ N_BI_c_467_n N_BI_c_506_p N_BI_c_479_n Vss PM_G5_XOR3_N1_BI
x_PM_G5_XOR3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_532_n
+ N_AI_c_566_p N_AI_c_522_n N_AI_c_523_n N_AI_c_537_n N_AI_c_527_n N_AI_c_528_n
+ N_AI_c_529_n N_AI_c_540_n Vss PM_G5_XOR3_N1_AI
x_PM_G5_XOR3_N1_B N_B_XI5.X0_CG N_B_XI6.X0_CG N_B_XI4.X0_CG N_B_XI3.X0_CG
+ N_B_c_576_n N_B_c_578_n N_B_c_590_n N_B_c_648_n N_B_c_611_n N_B_c_579_n B
+ N_B_c_615_n N_B_c_583_n N_B_c_580_n N_B_c_620_n N_B_c_621_n N_B_c_581_n
+ N_B_c_602_n N_B_c_603_n N_B_c_585_n N_B_c_645_n N_B_c_586_n Vss
+ PM_G5_XOR3_N1_B
x_PM_G5_XOR3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_669_n Z Vss PM_G5_XOR3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_C_XI9.X0_CG 9.6041e-19
cc_2 N_VDD_c_2_p N_C_XI9.X0_CG 8.03148e-19
cc_3 N_VDD_XI9.X0_PGD N_C_c_127_n 4.16623e-19
cc_4 N_VDD_c_4_p N_C_c_127_n 9.6041e-19
cc_5 N_VDD_c_5_p N_C_c_127_n 0.00125128f
cc_6 N_VDD_c_6_p C 4.36744e-19
cc_7 N_VDD_c_5_p C 0.00161703f
cc_8 N_VDD_c_6_p N_C_c_132_n 3.66936e-19
cc_9 N_VDD_c_5_p N_C_c_132_n 2.84956e-19
cc_10 N_VDD_XI6.X0_S N_C_c_134_n 3.43419e-19
cc_11 N_VDD_c_11_p N_C_c_135_n 4.67477e-19
cc_12 N_VDD_c_12_p N_C_c_135_n 7.7658e-19
cc_13 N_VDD_XI9.X0_PGD N_VSS_XI10.X0_PGD 0.00173038f
cc_14 N_VDD_c_5_p N_VSS_XI9.X0_S 3.7884e-19
cc_15 N_VDD_XI5.X0_PGD N_VSS_XI8.X0_PGD 2.27468e-19
cc_16 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172148f
cc_17 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017188f
cc_18 N_VDD_XI7.X0_PGD N_VSS_XI6.X0_PGD 2.1536e-19
cc_19 N_VDD_c_19_p N_VSS_XI7.X0_S 4.04413e-19
cc_20 N_VDD_c_20_p N_VSS_c_191_n 0.00173038f
cc_21 N_VDD_c_21_p N_VSS_c_192_n 0.00172148f
cc_22 N_VDD_c_22_p N_VSS_c_192_n 2.51785e-19
cc_23 N_VDD_c_22_p N_VSS_c_194_n 3.71017e-19
cc_24 N_VDD_c_12_p N_VSS_c_195_n 2.35445e-19
cc_25 N_VDD_c_25_p N_VSS_c_196_n 0.0017188f
cc_26 N_VDD_c_26_p N_VSS_c_196_n 2.74208e-19
cc_27 N_VDD_c_27_p N_VSS_c_198_n 4.32468e-19
cc_28 N_VDD_c_5_p N_VSS_c_198_n 4.60511e-19
cc_29 N_VDD_c_29_p N_VSS_c_198_n 0.00130521f
cc_30 N_VDD_c_30_p N_VSS_c_198_n 4.5978e-19
cc_31 N_VDD_c_31_p N_VSS_c_198_n 3.98949e-19
cc_32 N_VDD_c_2_p N_VSS_c_198_n 3.48267e-19
cc_33 N_VDD_c_5_p N_VSS_c_204_n 4.58491e-19
cc_34 N_VDD_c_34_p N_VSS_c_204_n 2.25587e-19
cc_35 N_VDD_c_11_p N_VSS_c_204_n 7.77634e-19
cc_36 N_VDD_c_12_p N_VSS_c_204_n 3.28649e-19
cc_37 N_VDD_c_37_p N_VSS_c_208_n 4.0876e-19
cc_38 N_VDD_c_22_p N_VSS_c_208_n 0.00141228f
cc_39 N_VDD_c_39_p N_VSS_c_208_n 8.73606e-19
cc_40 N_VDD_c_40_p N_VSS_c_208_n 3.48267e-19
cc_41 N_VDD_c_11_p N_VSS_c_212_n 6.87451e-19
cc_42 N_VDD_c_26_p N_VSS_c_212_n 0.00141228f
cc_43 N_VDD_c_12_p N_VSS_c_212_n 0.00254823f
cc_44 N_VDD_c_44_p N_VSS_c_212_n 3.48267e-19
cc_45 N_VDD_c_39_p N_VSS_c_216_n 7.30795e-19
cc_46 N_VDD_c_19_p N_VSS_c_216_n 5.00098e-19
cc_47 N_VDD_c_27_p N_VSS_c_218_n 4.41003e-19
cc_48 N_VDD_c_31_p N_VSS_c_218_n 3.89161e-19
cc_49 N_VDD_c_2_p N_VSS_c_218_n 7.99831e-19
cc_50 N_VDD_c_37_p N_VSS_c_221_n 3.48267e-19
cc_51 N_VDD_c_22_p N_VSS_c_221_n 0.00112249f
cc_52 N_VDD_c_39_p N_VSS_c_221_n 3.99794e-19
cc_53 N_VDD_c_40_p N_VSS_c_221_n 8.07559e-19
cc_54 N_VDD_c_11_p N_VSS_c_225_n 3.82294e-19
cc_55 N_VDD_c_26_p N_VSS_c_225_n 0.00112249f
cc_56 N_VDD_c_12_p N_VSS_c_225_n 9.55109e-19
cc_57 N_VDD_c_44_p N_VSS_c_225_n 8.01441e-19
cc_58 N_VDD_c_6_p N_VSS_c_229_n 0.003116f
cc_59 N_VDD_c_27_p N_VSS_c_229_n 7.60301e-19
cc_60 N_VDD_c_60_p N_VSS_c_229_n 0.0010705f
cc_61 N_VDD_c_27_p N_VSS_c_232_n 0.00754268f
cc_62 N_VDD_c_31_p N_VSS_c_232_n 9.72927e-19
cc_63 N_VDD_c_5_p N_VSS_c_234_n 0.00967241f
cc_64 N_VDD_c_64_p N_VSS_c_235_n 0.00107121f
cc_65 N_VDD_c_30_p N_VSS_c_236_n 0.0081111f
cc_66 N_VDD_c_34_p N_VSS_c_236_n 7.52646e-19
cc_67 N_VDD_c_22_p N_VSS_c_236_n 0.00375883f
cc_68 N_VDD_c_68_p N_VSS_c_236_n 0.0014027f
cc_69 N_VDD_c_27_p N_VSS_c_240_n 0.00107333f
cc_70 N_VDD_c_5_p N_VSS_c_241_n 0.00142828f
cc_71 N_VDD_c_26_p N_VSS_c_241_n 0.00543165f
cc_72 N_VDD_c_72_p N_VSS_c_241_n 0.00106247f
cc_73 N_VDD_c_22_p N_VSS_c_244_n 0.00372698f
cc_74 N_VDD_c_19_p N_VSS_c_244_n 0.00347642f
cc_75 N_VDD_c_27_p N_VSS_c_246_n 0.00112682f
cc_76 N_VDD_c_5_p N_VSS_c_247_n 0.00104966f
cc_77 N_VDD_c_22_p N_VSS_c_248_n 7.74609e-19
cc_78 N_VDD_XI10.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_79 N_VDD_c_29_p N_CI_XI10.X0_D 3.72199e-19
cc_80 N_VDD_XI10.X0_S N_CI_c_317_n 3.48267e-19
cc_81 N_VDD_c_5_p N_CI_c_317_n 5.01863e-19
cc_82 N_VDD_c_29_p N_CI_c_317_n 5.226e-19
cc_83 N_VDD_c_31_p N_CI_c_317_n 4.13481e-19
cc_84 N_VDD_c_31_p N_CI_c_321_n 7.11597e-19
cc_85 N_VDD_c_34_p N_CI_c_321_n 7.78475e-19
cc_86 N_VDD_c_40_p N_A_XI7.X0_CG 0.00119068f
cc_87 N_VDD_XI7.X0_PGD N_A_c_378_n 3.90714e-19
cc_88 N_VDD_XI6.X0_S N_A_c_379_n 2.96819e-19
cc_89 N_VDD_XI7.X0_PGD N_A_c_379_n 2.39692e-19
cc_90 N_VDD_c_22_p N_A_c_379_n 5.16693e-19
cc_91 N_VDD_c_26_p N_A_c_379_n 4.57585e-19
cc_92 N_VDD_c_39_p N_A_c_379_n 5.97577e-19
cc_93 N_VDD_c_12_p N_A_c_379_n 4.47961e-19
cc_94 N_VDD_c_19_p N_A_c_379_n 4.69788e-19
cc_95 N_VDD_c_40_p N_A_c_379_n 4.46731e-19
cc_96 N_VDD_XI6.X0_S N_A_c_387_n 9.18655e-19
cc_97 N_VDD_c_12_p N_A_c_388_n 0.00610545f
cc_98 N_VDD_c_31_p N_A_c_389_n 8.33062e-19
cc_99 N_VDD_c_31_p N_A_c_390_n 6.30148e-19
cc_100 N_VDD_c_44_p N_A_c_390_n 5.39283e-19
cc_101 N_VDD_XI6.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_102 N_VDD_c_12_p N_BI_XI5.X0_D 3.48267e-19
cc_103 N_VDD_XI6.X0_S N_BI_c_460_n 3.48267e-19
cc_104 N_VDD_c_26_p N_BI_c_460_n 4.87462e-19
cc_105 N_VDD_c_12_p N_BI_c_460_n 5.0516e-19
cc_106 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_107 N_VDD_c_22_p N_AI_XI8.X0_D 4.04413e-19
cc_108 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.98495e-19
cc_109 N_VDD_c_109_p N_AI_c_522_n 2.98495e-19
cc_110 N_VDD_XI8.X0_S N_AI_c_523_n 3.48267e-19
cc_111 N_VDD_c_34_p N_AI_c_523_n 4.96286e-19
cc_112 N_VDD_c_22_p N_AI_c_523_n 4.84258e-19
cc_113 N_VDD_c_39_p N_AI_c_523_n 5.74209e-19
cc_114 N_VDD_c_39_p N_AI_c_527_n 2.15672e-19
cc_115 N_VDD_c_19_p N_AI_c_528_n 3.25291e-19
cc_116 N_VDD_c_22_p N_AI_c_529_n 2.81017e-19
cc_117 N_VDD_XI9.X0_PGD N_B_XI5.X0_CG 9.57243e-19
cc_118 N_VDD_c_44_p N_B_XI5.X0_CG 9.74645e-19
cc_119 N_VDD_XI5.X0_PGD N_B_c_576_n 3.9688e-19
cc_120 N_VDD_XI7.X0_PGD N_B_c_576_n 2.07132e-19
cc_121 N_VDD_c_121_p N_B_c_578_n 9.57243e-19
cc_122 N_VDD_c_31_p N_B_c_579_n 6.08224e-19
cc_123 N_VDD_c_40_p N_B_c_580_n 3.47237e-19
cc_124 N_VDD_c_12_p N_B_c_581_n 2.72308e-19
cc_125 N_C_c_127_n N_VSS_XI10.X0_PGD 4.16623e-19
cc_126 N_C_c_132_n N_VSS_c_250_n 6.87259e-19
cc_127 C N_VSS_c_198_n 4.80408e-19
cc_128 N_C_c_140_p N_VSS_c_198_n 3.9981e-19
cc_129 N_C_c_141_p N_VSS_c_198_n 2.54015e-19
cc_130 N_C_c_135_n N_VSS_c_204_n 0.00185659f
cc_131 N_C_c_135_n N_VSS_c_212_n 0.00161389f
cc_132 N_C_c_144_p N_VSS_c_218_n 0.0041277f
cc_133 C N_VSS_c_218_n 4.20453e-19
cc_134 N_C_c_132_n N_VSS_c_218_n 0.00184261f
cc_135 N_C_c_140_p N_VSS_c_229_n 4.01014e-19
cc_136 N_C_c_141_p N_VSS_c_229_n 2.65147e-19
cc_137 C N_VSS_c_234_n 3.52403e-19
cc_138 N_C_c_140_p N_VSS_c_234_n 0.00136475f
cc_139 N_C_c_135_n N_VSS_c_234_n 0.00239048f
cc_140 N_C_c_141_p N_VSS_c_234_n 5.40072e-19
cc_141 N_C_c_135_n N_VSS_c_241_n 0.00182168f
cc_142 N_C_c_135_n N_CI_c_317_n 0.00135409f
cc_143 N_C_c_135_n N_CI_c_321_n 0.0042263f
cc_144 N_C_c_156_p N_CI_c_325_n 6.92841e-19
cc_145 N_C_c_157_p N_A_c_387_n 0.00149093f
cc_146 N_C_c_134_n N_A_c_387_n 8.20481e-19
cc_147 N_C_c_135_n N_A_c_387_n 2.83242e-19
cc_148 N_C_c_160_p N_A_c_387_n 2.26175e-19
cc_149 N_C_c_157_p N_A_c_396_n 0.00194268f
cc_150 N_C_c_134_n N_A_c_396_n 9.18655e-19
cc_151 N_C_c_135_n N_A_c_396_n 4.77334e-19
cc_152 N_C_c_156_p N_A_c_396_n 0.00211066f
cc_153 N_C_c_160_p N_A_c_396_n 6.30333e-19
cc_154 N_C_c_156_p N_A_c_401_n 5.46695e-19
cc_155 N_C_c_135_n N_BI_c_460_n 0.00227671f
cc_156 N_C_c_135_n N_BI_c_464_n 0.00490342f
cc_157 N_C_c_156_p N_BI_c_464_n 0.0015987f
cc_158 N_C_c_160_p N_BI_c_464_n 0.0013513f
cc_159 N_C_c_156_p N_BI_c_467_n 9.86034e-19
cc_160 N_C_c_135_n N_B_c_579_n 2.53746e-19
cc_161 N_C_c_156_p N_B_c_583_n 2.11999e-19
cc_162 N_C_c_157_p N_B_c_581_n 4.78342e-19
cc_163 N_C_c_156_p N_B_c_585_n 5.08651e-19
cc_164 N_C_c_156_p N_B_c_586_n 0.00239488f
cc_165 N_C_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_166 N_C_c_157_p N_Z_XI2.X0_D 3.48267e-19
cc_167 N_C_c_179_p N_Z_XI2.X0_D 3.48267e-19
cc_168 N_C_c_134_n N_Z_XI2.X0_D 3.43419e-19
cc_169 N_C_XI3.X0_S N_Z_c_669_n 3.48267e-19
cc_170 N_C_c_157_p N_Z_c_669_n 3.23828e-19
cc_171 N_C_c_179_p N_Z_c_669_n 5.71075e-19
cc_172 N_VSS_XI9.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_173 N_VSS_c_204_n N_CI_XI10.X0_D 3.48267e-19
cc_174 N_VSS_XI7.X0_S N_CI_XI4.X0_S 3.43419e-19
cc_175 N_VSS_c_216_n N_CI_XI4.X0_S 3.48267e-19
cc_176 N_VSS_c_198_n N_CI_c_317_n 5.88914e-19
cc_177 N_VSS_c_204_n N_CI_c_317_n 8.48865e-19
cc_178 N_VSS_c_234_n N_CI_c_317_n 3.32126e-19
cc_179 N_VSS_XI7.X0_S N_CI_c_333_n 3.48267e-19
cc_180 N_VSS_c_216_n N_CI_c_333_n 7.99744e-19
cc_181 N_VSS_c_208_n N_CI_c_321_n 3.41088e-19
cc_182 N_VSS_c_244_n N_CI_c_321_n 4.44969e-19
cc_183 N_VSS_c_232_n N_CI_c_337_n 2.78598e-19
cc_184 N_VSS_c_236_n N_CI_c_337_n 0.00159458f
cc_185 N_VSS_c_216_n N_CI_c_339_n 0.00104291f
cc_186 N_VSS_c_221_n N_A_c_402_n 0.00297797f
cc_187 N_VSS_XI8.X0_PGD N_A_c_378_n 3.85826e-19
cc_188 N_VSS_XI7.X0_S N_A_c_379_n 9.18655e-19
cc_189 N_VSS_c_216_n N_A_c_379_n 0.00131738f
cc_190 N_VSS_c_241_n N_A_c_379_n 3.01443e-19
cc_191 N_VSS_c_244_n N_A_c_379_n 5.02211e-19
cc_192 N_VSS_c_208_n N_A_c_389_n 5.62647e-19
cc_193 N_VSS_c_221_n N_A_c_389_n 4.60973e-19
cc_194 N_VSS_c_288_p N_A_c_390_n 9.36847e-19
cc_195 N_VSS_c_208_n N_A_c_390_n 4.56568e-19
cc_196 N_VSS_c_221_n N_A_c_390_n 8.15819e-19
cc_197 N_VSS_XI9.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_198 N_VSS_XI9.X0_S N_BI_c_460_n 3.48267e-19
cc_199 N_VSS_c_204_n N_BI_c_460_n 7.98486e-19
cc_200 N_VSS_c_241_n N_BI_c_460_n 3.20743e-19
cc_201 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_202 N_VSS_XI6.X0_PGD N_AI_XI2.X0_PGD 2.8463e-19
cc_203 N_VSS_c_195_n N_AI_c_532_n 2.8463e-19
cc_204 N_VSS_XI7.X0_S N_AI_c_523_n 3.48267e-19
cc_205 N_VSS_c_208_n N_AI_c_523_n 0.00108072f
cc_206 N_VSS_c_216_n N_AI_c_523_n 0.00193557f
cc_207 N_VSS_c_244_n N_AI_c_523_n 3.6914e-19
cc_208 N_VSS_c_216_n N_AI_c_537_n 8.20606e-19
cc_209 N_VSS_c_244_n N_AI_c_528_n 9.54335e-19
cc_210 N_VSS_c_244_n N_AI_c_529_n 0.00515467f
cc_211 N_VSS_c_244_n N_AI_c_540_n 0.00185629f
cc_212 N_VSS_c_225_n N_B_XI6.X0_CG 0.00272012f
cc_213 N_VSS_XI8.X0_PGD N_B_c_576_n 2.07132e-19
cc_214 N_VSS_XI6.X0_PGD N_B_c_576_n 3.923e-19
cc_215 N_VSS_c_225_n N_B_c_590_n 0.00130195f
cc_216 N_VSS_c_212_n N_B_c_579_n 7.62066e-19
cc_217 N_VSS_c_212_n B 5.66975e-19
cc_218 N_VSS_c_225_n B 4.56568e-19
cc_219 N_VSS_c_225_n N_B_c_580_n 6.1245e-19
cc_220 N_VSS_c_216_n N_B_c_581_n 6.79536e-19
cc_221 N_CI_c_339_n N_A_c_379_n 6.20926e-19
cc_222 N_CI_c_321_n N_A_c_389_n 0.00116415f
cc_223 N_CI_c_339_n N_A_c_389_n 2.08707e-19
cc_224 N_CI_c_317_n N_BI_c_460_n 5.94242e-19
cc_225 N_CI_c_321_n N_BI_c_460_n 0.00302092f
cc_226 N_CI_c_333_n N_BI_c_464_n 3.50977e-19
cc_227 N_CI_c_321_n N_BI_c_464_n 0.00752744f
cc_228 N_CI_c_347_p N_BI_c_464_n 4.80593e-19
cc_229 N_CI_c_325_n N_BI_c_464_n 5.67893e-19
cc_230 N_CI_c_325_n N_BI_c_478_n 0.00102574f
cc_231 N_CI_c_325_n N_BI_c_479_n 2.55507e-19
cc_232 N_CI_c_321_n N_AI_c_523_n 8.44506e-19
cc_233 N_CI_c_339_n N_AI_c_523_n 0.00100365f
cc_234 N_CI_c_325_n N_AI_c_537_n 0.00169084f
cc_235 N_CI_c_333_n N_AI_c_528_n 8.33462e-19
cc_236 N_CI_c_347_p N_AI_c_528_n 7.14401e-19
cc_237 N_CI_c_356_p N_AI_c_528_n 2.16882e-19
cc_238 N_CI_c_325_n N_AI_c_528_n 5.16616e-19
cc_239 N_CI_c_321_n N_AI_c_529_n 0.00115159f
cc_240 N_CI_c_356_p N_AI_c_529_n 0.00241787f
cc_241 N_CI_c_317_n N_B_c_579_n 2.7112e-19
cc_242 N_CI_c_325_n N_B_c_583_n 7.18914e-19
cc_243 N_CI_c_333_n N_B_c_581_n 8.80932e-19
cc_244 N_CI_c_321_n N_B_c_581_n 0.00348609f
cc_245 N_CI_c_347_p N_B_c_581_n 2.27019e-19
cc_246 N_CI_c_325_n N_B_c_581_n 2.27123e-19
cc_247 N_CI_c_321_n N_B_c_602_n 0.00142048f
cc_248 N_CI_c_339_n N_B_c_603_n 3.62522e-19
cc_249 N_CI_c_339_n N_B_c_585_n 4.56062e-19
cc_250 N_CI_c_325_n N_B_c_585_n 0.00270237f
cc_251 N_CI_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_252 N_CI_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_253 N_CI_c_333_n N_Z_XI4.X0_D 3.48267e-19
cc_254 N_CI_c_373_p N_Z_XI4.X0_D 3.48267e-19
cc_255 N_CI_XI4.X0_S N_Z_c_669_n 3.48267e-19
cc_256 N_CI_c_333_n N_Z_c_669_n 5.68744e-19
cc_257 N_CI_c_373_p N_Z_c_669_n 6.06579e-19
cc_258 N_A_c_396_n N_BI_c_480_n 3.17089e-19
cc_259 N_A_XI3.X0_PGD N_BI_c_481_n 8.79767e-19
cc_260 N_A_c_379_n N_BI_c_460_n 4.32688e-19
cc_261 N_A_c_387_n N_BI_c_464_n 9.32646e-19
cc_262 N_A_c_396_n N_BI_c_464_n 5.00869e-19
cc_263 N_A_c_396_n N_BI_c_478_n 3.33012e-19
cc_264 N_A_c_387_n N_BI_c_486_n 3.37713e-19
cc_265 N_A_XI3.X0_PGD N_BI_c_487_n 0.00133285f
cc_266 N_A_c_396_n N_BI_c_467_n 0.00106538f
cc_267 N_A_c_379_n N_AI_XI8.X0_D 9.18655e-19
cc_268 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174819f
cc_269 N_A_c_387_n N_AI_XI2.X0_PGD 8.52417e-19
cc_270 N_A_c_428_p N_AI_c_532_n 0.00199595f
cc_271 N_A_c_396_n N_AI_c_532_n 0.00123184f
cc_272 N_A_c_430_p N_AI_c_522_n 0.00202022f
cc_273 N_A_c_379_n N_AI_c_523_n 0.00136181f
cc_274 N_A_c_379_n N_AI_c_529_n 2.67536e-19
cc_275 N_A_XI3.X0_PGD N_B_XI3.X0_CG 8.79767e-19
cc_276 N_A_c_434_p N_B_XI3.X0_CG 0.00237738f
cc_277 N_A_c_378_n N_B_c_576_n 0.0036024f
cc_278 N_A_c_379_n N_B_c_576_n 5.40888e-19
cc_279 N_A_c_390_n N_B_c_578_n 4.08399e-19
cc_280 N_A_c_434_p N_B_c_611_n 0.00115102f
cc_281 N_A_c_387_n N_B_c_579_n 6.16253e-19
cc_282 N_A_c_379_n B 7.07944e-19
cc_283 N_A_c_387_n B 5.00495e-19
cc_284 N_A_c_379_n N_B_c_615_n 2.41829e-19
cc_285 N_A_c_401_n N_B_c_583_n 8.44727e-19
cc_286 N_A_c_434_p N_B_c_583_n 4.84491e-19
cc_287 N_A_c_378_n N_B_c_580_n 2.87365e-19
cc_288 N_A_c_387_n N_B_c_580_n 6.85754e-19
cc_289 N_A_c_379_n N_B_c_620_n 3.8563e-19
cc_290 N_A_XI3.X0_PGD N_B_c_621_n 0.00133285f
cc_291 N_A_c_401_n N_B_c_621_n 4.67029e-19
cc_292 N_A_c_434_p N_B_c_621_n 0.0014909f
cc_293 N_A_c_387_n N_B_c_581_n 0.00225059f
cc_294 N_A_c_396_n N_B_c_581_n 8.88958e-19
cc_295 N_A_c_379_n N_B_c_602_n 0.00244205f
cc_296 N_A_c_396_n N_Z_XI2.X0_D 6.94686e-19
cc_297 N_A_XI3.X0_PGD N_Z_c_669_n 6.30408e-19
cc_298 N_A_c_387_n N_Z_c_669_n 0.00124827f
cc_299 N_A_c_396_n N_Z_c_669_n 0.00121415f
cc_300 N_BI_XI2.X0_CG N_AI_XI2.X0_PGD 8.63152e-19
cc_301 N_BI_c_486_n N_AI_XI2.X0_PGD 0.00133285f
cc_302 N_BI_c_464_n N_AI_c_529_n 3.64122e-19
cc_303 N_BI_c_464_n N_B_c_579_n 0.00139574f
cc_304 N_BI_c_464_n N_B_c_615_n 6.02887e-19
cc_305 N_BI_c_479_n N_B_c_615_n 3.05615e-19
cc_306 N_BI_c_478_n N_B_c_583_n 0.00178808f
cc_307 N_BI_c_467_n N_B_c_583_n 0.00156529f
cc_308 N_BI_c_464_n N_B_c_620_n 4.56568e-19
cc_309 N_BI_c_486_n N_B_c_620_n 0.00266354f
cc_310 N_BI_c_487_n N_B_c_620_n 7.16621e-19
cc_311 N_BI_c_478_n N_B_c_621_n 4.56568e-19
cc_312 N_BI_c_486_n N_B_c_621_n 6.17967e-19
cc_313 N_BI_c_487_n N_B_c_621_n 0.00243716f
cc_314 N_BI_c_464_n N_B_c_581_n 0.00427216f
cc_315 N_BI_c_464_n N_B_c_603_n 3.15526e-19
cc_316 N_BI_c_467_n N_B_c_603_n 0.00129112f
cc_317 N_BI_c_506_p N_B_c_603_n 0.0034245f
cc_318 N_BI_c_464_n N_B_c_585_n 4.99817e-19
cc_319 N_BI_c_467_n N_B_c_585_n 7.12768e-19
cc_320 N_BI_c_479_n N_B_c_585_n 7.15853e-19
cc_321 N_BI_c_506_p N_B_c_645_n 0.00229162f
cc_322 N_BI_c_464_n N_B_c_586_n 0.00139788f
cc_323 N_BI_c_467_n N_B_c_586_n 8.65145e-19
cc_324 N_BI_c_464_n N_Z_c_669_n 0.00138937f
cc_325 N_BI_c_478_n N_Z_c_669_n 0.00157561f
cc_326 N_BI_c_486_n N_Z_c_669_n 8.66889e-19
cc_327 N_BI_c_467_n N_Z_c_669_n 0.00100271f
cc_328 N_BI_c_506_p N_Z_c_669_n 0.00210866f
cc_329 N_BI_c_479_n N_Z_c_669_n 9.67357e-19
cc_330 N_AI_XI2.X0_PGD N_B_c_648_n 8.79767e-19
cc_331 N_AI_c_527_n N_B_c_648_n 0.00234569f
cc_332 N_AI_c_537_n N_B_c_615_n 5.49665e-19
cc_333 N_AI_c_527_n N_B_c_615_n 4.745e-19
cc_334 N_AI_XI2.X0_PGD N_B_c_620_n 0.00133285f
cc_335 N_AI_c_566_p N_B_c_620_n 7.60534e-19
cc_336 N_AI_c_537_n N_B_c_620_n 4.46045e-19
cc_337 N_AI_c_527_n N_B_c_620_n 0.00166302f
cc_338 N_AI_c_528_n N_B_c_581_n 0.00120142f
cc_339 N_AI_c_529_n N_B_c_581_n 3.28172e-19
cc_340 N_AI_c_529_n N_B_c_602_n 2.8335e-19
cc_341 N_AI_c_537_n N_B_c_603_n 4.27113e-19
cc_342 N_AI_XI2.X0_PGD N_Z_c_669_n 3.26804e-19
cc_343 N_B_c_615_n N_Z_c_669_n 0.0013937f
cc_344 N_B_c_583_n N_Z_c_669_n 0.00139745f
cc_345 N_B_c_620_n N_Z_c_669_n 8.66889e-19
cc_346 N_B_c_621_n N_Z_c_669_n 8.66889e-19
cc_347 N_B_c_603_n N_Z_c_669_n 4.72173e-19
*
.ends
*
*
.subckt XOR3_HPNW4 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XOR3_N1_2
.ends
*
* File: G3_AND2_N2.pex.netlist
* Created: Mon Feb 28 10:46:36 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_AND2_N2_VSS 2 3 5 6 8 9 11 13 27 28 30 49 62 67 73 78 83 88 97 102
+ 111 112 116 117 122 128 130 135 136 137 139 Vss
c70 137 Vss 3.78257e-19
c71 136 Vss 3.62111e-19
c72 135 Vss 0.00438377f
c73 130 Vss 0.00256681f
c74 128 Vss 0.00549491f
c75 122 Vss 0.00414054f
c76 117 Vss 8.38241e-19
c77 116 Vss 0.00175385f
c78 112 Vss 7.28672e-19
c79 111 Vss 0.00525523f
c80 102 Vss 0.00402938f
c81 97 Vss 0.00450731f
c82 88 Vss 7.10513e-22
c83 83 Vss 4.8239e-19
c84 78 Vss 0.00106653f
c85 73 Vss 0.00125808f
c86 67 Vss 0.00537538f
c87 62 Vss 0.00490594f
c88 58 Vss 0.0299355f
c89 57 Vss 0.0299355f
c90 50 Vss 0.0347118f
c91 49 Vss 0.0994217f
c92 41 Vss 0.106723f
c93 35 Vss 0.0688517f
c94 30 Vss 5.38535e-20
c95 28 Vss 0.0340588f
c96 27 Vss 0.064644f
c97 11 Vss 0.134525f
c98 9 Vss 0.134971f
c99 8 Vss 0.133544f
c100 6 Vss 0.134177f
c101 5 Vss 0.138048f
c102 3 Vss 0.135913f
r103 135 139 0.326018
r104 134 135 5.08479
r105 130 134 0.655813
r106 129 137 0.494161
r107 128 139 0.326018
r108 128 129 10.1279
r109 124 137 0.128424
r110 123 136 0.494161
r111 122 137 0.494161
r112 122 123 10.378
r113 118 136 0.128424
r114 116 136 0.494161
r115 116 117 4.33457
r116 111 117 0.652036
r117 110 112 0.655813
r118 110 111 16.6297
r119 88 130 1.82344
r120 83 102 1.16709
r121 83 124 2.66743
r122 78 97 1.16709
r123 78 118 2.16729
r124 73 112 1.82344
r125 67 88 1.16709
r126 62 73 1.16709
r127 52 102 0.0476429
r128 50 52 1.45875
r129 49 53 0.652036
r130 49 52 1.45875
r131 46 50 0.652036
r132 42 58 0.494161
r133 41 43 0.652036
r134 41 42 2.9175
r135 37 58 0.128424
r136 36 57 0.494161
r137 35 58 0.494161
r138 35 36 2.8008
r139 31 57 0.128424
r140 30 97 0.238214
r141 28 30 1.4004
r142 27 57 0.494161
r143 27 30 1.5171
r144 24 28 0.652036
r145 13 67 0.185659
r146 11 46 3.8511
r147 9 53 3.8511
r148 8 43 3.8511
r149 6 37 3.8511
r150 5 24 3.8511
r151 3 31 3.8511
r152 2 62 0.185659
.ends

.subckt PM_G3_AND2_N2_VDD 1 3 5 7 8 10 24 26 33 43 48 53 55 56 60 62 63 66 70 72
+ 74 76 78 79 81 87 96 Vss
c85 96 Vss 0.00462548f
c86 87 Vss 0.00521601f
c87 79 Vss 4.60053e-19
c88 78 Vss 4.52364e-19
c89 76 Vss 0.00122604f
c90 74 Vss 6.12561e-19
c91 72 Vss 0.00375739f
c92 70 Vss 0.001382f
c93 66 Vss 0.00251556f
c94 63 Vss 8.66752e-19
c95 62 Vss 0.00754689f
c96 60 Vss 0.0017718f
c97 57 Vss 0.00173794f
c98 56 Vss 0.010708f
c99 55 Vss 0.00235908f
c100 53 Vss 0.00679887f
c101 48 Vss 0.00711219f
c102 43 Vss 0.00386059f
c103 33 Vss 0.0357726f
c104 32 Vss 0.102409f
c105 26 Vss 0.170515f
c106 24 Vss 0.0339269f
c107 10 Vss 0.136393f
c108 8 Vss 0.13497f
c109 7 Vss 0.00143442f
c110 1 Vss 0.117228f
r111 76 96 1.16709
r112 74 81 0.326018
r113 74 76 2.66743
r114 73 79 0.494161
r115 72 81 0.326018
r116 72 73 7.46046
r117 68 79 0.128424
r118 68 70 5.75164
r119 66 87 1.16709
r120 64 66 3.83443
r121 62 79 0.494161
r122 62 63 13.0037
r123 58 78 0.0828784
r124 58 60 1.82344
r125 56 64 0.652036
r126 56 57 10.0862
r127 55 63 0.652036
r128 54 78 0.551426
r129 54 55 5.08479
r130 53 78 0.551426
r131 52 57 0.652036
r132 52 53 13.0454
r133 48 70 1.16709
r134 43 60 1.16709
r135 35 96 0.0476429
r136 33 35 1.45875
r137 32 36 0.652036
r138 32 35 1.45875
r139 28 33 0.652036
r140 26 87 0.428786
r141 24 26 5.3682
r142 20 24 0.652036
r143 10 36 3.8511
r144 8 28 3.8511
r145 7 48 0.185659
r146 5 48 0.185659
r147 3 43 0.185659
r148 1 20 3.1509
.ends

.subckt PM_G3_AND2_N2_A 2 4 10 13 18 21 26 31 Vss
c26 31 Vss 0.00351072f
c27 26 Vss 0.00323449f
c28 18 Vss 9.2489e-19
c29 13 Vss 0.112394f
c30 2 Vss 0.112081f
r31 23 31 1.16709
r32 21 23 2.95918
r33 18 26 1.16709
r34 18 21 2.41736
r35 13 31 0.50025
r36 10 26 0.50025
r37 4 13 3.09255
r38 2 10 3.09255
.ends

.subckt PM_G3_AND2_N2_NET1 2 4 6 8 10 24 27 38 42 46 50 52 56 68 Vss
c52 68 Vss 0.00584624f
c53 58 Vss 1.47786e-19
c54 56 Vss 0.00230674f
c55 52 Vss 0.00700301f
c56 50 Vss 0.00103961f
c57 46 Vss 7.16542e-19
c58 42 Vss 0.00585482f
c59 38 Vss 0.00349773f
c60 27 Vss 9.81095e-20
c61 24 Vss 0.227317f
c62 21 Vss 0.125908f
c63 19 Vss 0.0247918f
c64 10 Vss 0.139046f
c65 6 Vss 0.00143442f
r66 56 68 1.16709
r67 54 56 3.45932
r68 53 58 0.128424
r69 52 54 0.652036
r70 52 53 7.46046
r71 48 58 0.494161
r72 48 50 6.54354
r73 44 58 0.494161
r74 44 46 3.83443
r75 42 50 1.16709
r76 38 46 1.16709
r77 27 68 0.0476429
r78 25 27 0.326018
r79 25 27 0.1167
r80 24 28 0.652036
r81 24 27 6.7686
r82 21 68 0.357321
r83 19 27 0.326018
r84 19 21 0.40845
r85 10 28 3.8511
r86 8 21 3.44265
r87 6 42 0.185659
r88 4 42 0.185659
r89 2 38 0.185659
.ends

.subckt PM_G3_AND2_N2_B 2 4 10 11 14 21 Vss
c26 21 Vss 3.50736e-19
c27 14 Vss 0.181075f
c28 11 Vss 0.0348746f
c29 10 Vss 0.288064f
c30 2 Vss 0.277377f
r31 18 21 0.0729375
r32 14 18 1.16709
r33 12 14 2.1006
r34 10 12 0.652036
r35 10 11 8.92755
r36 7 11 0.652036
r37 4 14 4.3179
r38 2 7 8.57745
.ends

.subckt PM_G3_AND2_N2_Z 2 4 13 18 Vss
c13 13 Vss 0.0052353f
c14 4 Vss 0.00143442f
r15 13 18 1.16709
r16 4 13 0.185659
r17 2 13 0.185659
.ends

.subckt G3_AND2_N2  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI5.X0 N_NET1_XI5.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_B_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW8
XI10.X0 N_NET1_XI10.X0_D N_VSS_XI10.X0_PGD N_A_XI10.X0_CG N_VSS_XI10.X0_PGS
+ N_VDD_XI10.X0_S TIGFET_HPNW8
XI6.X0 N_NET1_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGS
+ N_VDD_XI6.X0_S TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VSS_XI4.X0_PGD N_NET1_XI4.X0_CG N_VSS_XI4.X0_PGS
+ N_VDD_XI4.X0_S TIGFET_HPNW8
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_NET1_XI3.X0_CG N_VDD_XI3.X0_PGS
+ N_VSS_XI3.X0_S TIGFET_HPNW8
*
x_PM_G3_AND2_N2_VSS N_VSS_XI5.X0_S N_VSS_XI10.X0_PGD N_VSS_XI10.X0_PGS
+ N_VSS_XI6.X0_PGD N_VSS_XI6.X0_PGS N_VSS_XI4.X0_PGD N_VSS_XI4.X0_PGS
+ N_VSS_XI3.X0_S N_VSS_c_13_p N_VSS_c_14_p N_VSS_c_46_p N_VSS_c_2_p N_VSS_c_3_p
+ N_VSS_c_65_p N_VSS_c_4_p N_VSS_c_8_p N_VSS_c_24_p N_VSS_c_66_p N_VSS_c_9_p
+ N_VSS_c_26_p N_VSS_c_5_p N_VSS_c_6_p N_VSS_c_17_p N_VSS_c_20_p N_VSS_c_18_p
+ N_VSS_c_32_p N_VSS_c_70_p N_VSS_c_37_p N_VSS_c_19_p N_VSS_c_33_p VSS Vss
+ PM_G3_AND2_N2_VSS
x_PM_G3_AND2_N2_VDD N_VDD_XI5.X0_PGD N_VDD_XI10.X0_S N_VDD_XI6.X0_S
+ N_VDD_XI4.X0_S N_VDD_XI3.X0_PGD N_VDD_XI3.X0_PGS N_VDD_c_148_p N_VDD_c_130_p
+ N_VDD_c_72_n N_VDD_c_125_p N_VDD_c_126_p N_VDD_c_73_n N_VDD_c_77_n
+ N_VDD_c_81_n N_VDD_c_82_n N_VDD_c_83_n N_VDD_c_90_n N_VDD_c_123_p N_VDD_c_91_n
+ N_VDD_c_98_n N_VDD_c_104_n N_VDD_c_105_n N_VDD_c_108_n N_VDD_c_109_n VDD
+ N_VDD_c_119_p N_VDD_c_110_n Vss PM_G3_AND2_N2_VDD
x_PM_G3_AND2_N2_A N_A_XI5.X0_CG N_A_XI10.X0_CG N_A_c_164_n N_A_c_156_n
+ N_A_c_157_n A N_A_c_167_n N_A_c_160_n Vss PM_G3_AND2_N2_A
x_PM_G3_AND2_N2_NET1 N_NET1_XI5.X0_D N_NET1_XI10.X0_D N_NET1_XI6.X0_D
+ N_NET1_XI4.X0_CG N_NET1_XI3.X0_CG N_NET1_c_182_n N_NET1_c_183_n N_NET1_c_184_n
+ N_NET1_c_199_n N_NET1_c_186_n N_NET1_c_189_n N_NET1_c_190_n N_NET1_c_191_n
+ N_NET1_c_193_n Vss PM_G3_AND2_N2_NET1
x_PM_G3_AND2_N2_B N_B_XI5.X0_PGS N_B_XI6.X0_CG N_B_c_234_n N_B_c_236_n
+ N_B_c_241_n B Vss PM_G3_AND2_N2_B
x_PM_G3_AND2_N2_Z N_Z_XI4.X0_D N_Z_XI3.X0_D N_Z_c_260_n Z Vss PM_G3_AND2_N2_Z
cc_1 N_VSS_XI4.X0_PGD N_VDD_XI3.X0_PGD 0.00195824f
cc_2 N_VSS_c_2_p N_VDD_c_72_n 0.00195824f
cc_3 N_VSS_c_3_p N_VDD_c_73_n 9.5668e-19
cc_4 N_VSS_c_4_p N_VDD_c_73_n 0.00165395f
cc_5 N_VSS_c_5_p N_VDD_c_73_n 0.00670587f
cc_6 N_VSS_c_6_p N_VDD_c_73_n 0.00189531f
cc_7 N_VSS_XI10.X0_PGS N_VDD_c_77_n 2.75457e-19
cc_8 N_VSS_c_8_p N_VDD_c_77_n 4.50283e-19
cc_9 N_VSS_c_9_p N_VDD_c_77_n 3.70842e-19
cc_10 N_VSS_c_5_p N_VDD_c_77_n 0.00345577f
cc_11 N_VSS_c_4_p N_VDD_c_81_n 0.00247496f
cc_12 N_VSS_c_4_p N_VDD_c_82_n 4.32396e-19
cc_13 N_VSS_c_13_p N_VDD_c_83_n 0.00151774f
cc_14 N_VSS_c_14_p N_VDD_c_83_n 3.51214e-19
cc_15 N_VSS_c_8_p N_VDD_c_83_n 0.00161703f
cc_16 N_VSS_c_9_p N_VDD_c_83_n 2.03837e-19
cc_17 N_VSS_c_17_p N_VDD_c_83_n 0.00348097f
cc_18 N_VSS_c_18_p N_VDD_c_83_n 0.0059139f
cc_19 N_VSS_c_19_p N_VDD_c_83_n 7.61747e-19
cc_20 N_VSS_c_20_p N_VDD_c_90_n 0.00107346f
cc_21 N_VSS_XI6.X0_PGS N_VDD_c_91_n 2.23834e-19
cc_22 N_VSS_XI4.X0_PGS N_VDD_c_91_n 2.29703e-19
cc_23 N_VSS_c_8_p N_VDD_c_91_n 6.50938e-19
cc_24 N_VSS_c_24_p N_VDD_c_91_n 0.00193467f
cc_25 N_VSS_c_9_p N_VDD_c_91_n 2.56577e-19
cc_26 N_VSS_c_26_p N_VDD_c_91_n 9.55109e-19
cc_27 N_VSS_c_5_p N_VDD_c_91_n 3.54686e-19
cc_28 N_VSS_c_2_p N_VDD_c_98_n 4.82224e-19
cc_29 N_VSS_c_24_p N_VDD_c_98_n 0.00118142f
cc_30 N_VSS_c_26_p N_VDD_c_98_n 2.13453e-19
cc_31 N_VSS_c_18_p N_VDD_c_98_n 0.00133442f
cc_32 N_VSS_c_32_p N_VDD_c_98_n 0.00433318f
cc_33 N_VSS_c_33_p N_VDD_c_98_n 8.13487e-19
cc_34 N_VSS_c_32_p N_VDD_c_104_n 0.00157826f
cc_35 N_VSS_c_24_p N_VDD_c_105_n 9.21598e-19
cc_36 N_VSS_c_26_p N_VDD_c_105_n 3.82294e-19
cc_37 N_VSS_c_37_p N_VDD_c_105_n 5.22507e-19
cc_38 N_VSS_c_5_p N_VDD_c_108_n 0.00100712f
cc_39 N_VSS_c_18_p N_VDD_c_109_n 9.86755e-19
cc_40 N_VSS_c_24_p N_VDD_c_110_n 3.48267e-19
cc_41 N_VSS_c_26_p N_VDD_c_110_n 6.46219e-19
cc_42 N_VSS_c_9_p N_A_c_156_n 0.00249847f
cc_43 N_VSS_c_8_p N_A_c_157_n 2.94885e-19
cc_44 N_VSS_c_9_p N_A_c_157_n 3.71222e-19
cc_45 N_VSS_c_5_p N_A_c_157_n 0.00147463f
cc_46 N_VSS_c_46_p N_A_c_160_n 3.96531e-19
cc_47 N_VSS_c_8_p N_A_c_160_n 2.87758e-19
cc_48 N_VSS_c_9_p N_A_c_160_n 8.98435e-19
cc_49 N_VSS_XI4.X0_PGD N_NET1_c_182_n 4.26252e-19
cc_50 N_VSS_c_26_p N_NET1_c_183_n 9.4551e-19
cc_51 N_VSS_c_3_p N_NET1_c_184_n 3.43419e-19
cc_52 N_VSS_c_4_p N_NET1_c_184_n 3.48267e-19
cc_53 N_VSS_c_3_p N_NET1_c_186_n 3.48267e-19
cc_54 N_VSS_c_4_p N_NET1_c_186_n 8.50248e-19
cc_55 N_VSS_c_5_p N_NET1_c_186_n 5.59972e-19
cc_56 N_VSS_c_18_p N_NET1_c_189_n 2.3523e-19
cc_57 N_VSS_c_18_p N_NET1_c_190_n 4.47676e-19
cc_58 N_VSS_c_24_p N_NET1_c_191_n 5.58211e-19
cc_59 N_VSS_c_26_p N_NET1_c_191_n 3.49408e-19
cc_60 N_VSS_c_24_p N_NET1_c_193_n 3.2351e-19
cc_61 N_VSS_c_26_p N_NET1_c_193_n 2.68747e-19
cc_62 N_VSS_XI10.X0_PGD N_B_c_234_n 8.28117e-19
cc_63 N_VSS_XI6.X0_PGD N_B_c_234_n 8.28117e-19
cc_64 N_VSS_XI10.X0_PGS N_B_c_236_n 9.94582e-19
cc_65 N_VSS_c_65_p N_Z_c_260_n 3.43419e-19
cc_66 N_VSS_c_66_p N_Z_c_260_n 3.48267e-19
cc_67 N_VSS_c_65_p Z 3.48267e-19
cc_68 N_VSS_c_66_p Z 4.99861e-19
cc_69 N_VSS_c_32_p Z 2.34298e-19
cc_70 N_VSS_c_70_p Z 2.7826e-19
cc_71 N_VDD_XI5.X0_PGD N_A_XI5.X0_CG 5.26351e-19
cc_72 N_VDD_c_81_n N_A_c_164_n 3.14632e-19
cc_73 N_VDD_c_73_n N_A_c_157_n 0.00285022f
cc_74 N_VDD_c_81_n N_A_c_157_n 5.83159e-19
cc_75 N_VDD_XI5.X0_PGD N_A_c_167_n 2.78309e-19
cc_76 N_VDD_c_73_n N_A_c_167_n 3.66936e-19
cc_77 N_VDD_c_81_n N_A_c_167_n 3.4118e-19
cc_78 N_VDD_c_119_p N_A_c_167_n 4.44265e-19
cc_79 N_VDD_c_73_n N_A_c_160_n 4.70132e-19
cc_80 N_VDD_XI3.X0_PGD N_NET1_c_182_n 4.29017e-19
cc_81 N_VDD_c_81_n N_NET1_c_184_n 9.18655e-19
cc_82 N_VDD_c_123_p N_NET1_c_184_n 8.835e-19
cc_83 N_VDD_c_119_p N_NET1_c_184_n 0.00132057f
cc_84 N_VDD_c_125_p N_NET1_c_199_n 3.43419e-19
cc_85 N_VDD_c_126_p N_NET1_c_199_n 3.43419e-19
cc_86 N_VDD_c_82_n N_NET1_c_199_n 3.72199e-19
cc_87 N_VDD_c_83_n N_NET1_c_199_n 3.02646e-19
cc_88 N_VDD_c_91_n N_NET1_c_199_n 3.48267e-19
cc_89 N_VDD_c_130_p N_NET1_c_186_n 7.85476e-19
cc_90 N_VDD_c_73_n N_NET1_c_186_n 9.00704e-19
cc_91 N_VDD_c_81_n N_NET1_c_186_n 0.00168791f
cc_92 N_VDD_c_123_p N_NET1_c_186_n 0.00355804f
cc_93 N_VDD_c_119_p N_NET1_c_186_n 8.835e-19
cc_94 N_VDD_c_125_p N_NET1_c_189_n 3.48267e-19
cc_95 N_VDD_c_126_p N_NET1_c_189_n 3.48267e-19
cc_96 N_VDD_c_82_n N_NET1_c_189_n 8.08807e-19
cc_97 N_VDD_c_83_n N_NET1_c_189_n 4.24175e-19
cc_98 N_VDD_c_91_n N_NET1_c_189_n 7.1497e-19
cc_99 N_VDD_c_130_p N_NET1_c_190_n 3.97408e-19
cc_100 N_VDD_c_126_p N_NET1_c_190_n 2.52932e-19
cc_101 N_VDD_c_123_p N_NET1_c_190_n 0.001476f
cc_102 N_VDD_c_91_n N_NET1_c_190_n 5.44012e-19
cc_103 N_VDD_c_119_p N_NET1_c_190_n 0.00114101f
cc_104 N_VDD_XI5.X0_PGD N_B_XI5.X0_PGS 0.00153355f
cc_105 N_VDD_c_73_n N_B_XI5.X0_PGS 7.45044e-19
cc_106 N_VDD_c_81_n N_B_XI5.X0_PGS 3.02077e-19
cc_107 N_VDD_c_148_p N_B_c_234_n 0.00419437f
cc_108 N_VDD_c_119_p N_B_c_241_n 7.17663e-19
cc_109 N_VDD_c_126_p N_Z_c_260_n 3.43419e-19
cc_110 N_VDD_c_91_n N_Z_c_260_n 3.48267e-19
cc_111 N_VDD_c_98_n N_Z_c_260_n 3.02646e-19
cc_112 N_VDD_c_126_p Z 3.48267e-19
cc_113 N_VDD_c_91_n Z 7.09569e-19
cc_114 N_VDD_c_98_n Z 4.04319e-19
cc_115 N_A_c_157_n N_NET1_c_186_n 0.00799902f
cc_116 N_A_c_167_n N_NET1_c_186_n 8.66889e-19
cc_117 N_A_c_160_n N_NET1_c_189_n 9.68342e-19
cc_118 N_A_XI5.X0_CG N_B_XI5.X0_PGS 4.87172e-19
cc_119 N_A_c_157_n N_B_XI5.X0_PGS 4.74011e-19
cc_120 N_A_c_167_n N_B_XI5.X0_PGS 5.6636e-19
cc_121 N_A_c_157_n N_B_c_234_n 2.0632e-19
cc_122 N_A_c_167_n N_B_c_234_n 7.2846e-19
cc_123 N_A_c_160_n N_B_c_234_n 0.00228839f
cc_124 N_A_c_160_n N_B_c_241_n 9.27569e-19
cc_125 N_NET1_c_199_n N_B_c_234_n 3.74089e-19
cc_126 N_NET1_c_189_n N_B_c_234_n 3.943e-19
cc_127 N_NET1_c_190_n N_B_c_234_n 2.82146e-19
cc_128 N_NET1_c_189_n N_B_c_241_n 0.00116203f
cc_129 N_NET1_c_190_n N_B_c_241_n 5.60175e-19
cc_130 N_NET1_c_191_n N_B_c_241_n 3.86148e-19
cc_131 N_NET1_c_193_n N_B_c_241_n 0.00196155f
cc_132 N_NET1_c_189_n B 0.00147455f
cc_133 N_NET1_c_190_n B 8.26881e-19
cc_134 N_NET1_c_191_n B 5.75904e-19
cc_135 N_NET1_c_193_n B 3.48267e-19
cc_136 N_NET1_c_182_n N_Z_c_260_n 6.55689e-19
*
.ends
*
*
.subckt AND2_HPNW8 A B Y VDD VSS
xgate (VSS VDD A B Y) G3_AND2_N2
.ends
*
* File: G2_AOI21_N2.pex.netlist
* Created: Mon Apr 11 18:40:10 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_AOI21_N2_VSS 2 4 6 8 19 30 35 38 43 48 57 66 67 69 77 78 79 84 86
+ 88 89 Vss
c51 89 Vss 4.28045e-19
c52 86 Vss 0.00486026f
c53 84 Vss 0.00155386f
c54 79 Vss 0.00128356f
c55 78 Vss 4.65637e-19
c56 77 Vss 0.00250049f
c57 69 Vss 0.00102564f
c58 67 Vss 0.00986383f
c59 66 Vss 0.00273179f
c60 65 Vss 0.00133186f
c61 57 Vss 0.00579208f
c62 48 Vss 2.73256e-19
c63 43 Vss 0.00178422f
c64 38 Vss 0.00142279f
c65 35 Vss 0.00389683f
c66 30 Vss 0.00549227f
c67 25 Vss 0.0828998f
c68 19 Vss 0.0350566f
c69 18 Vss 0.0688416f
c70 8 Vss 0.135691f
c71 4 Vss 0.134006f
r72 85 89 0.551426
r73 85 86 15.5878
r74 84 89 0.551426
r75 83 84 4.58464
r76 79 89 0.0828784
r77 77 86 0.652036
r78 77 78 4.33457
r79 73 78 0.652036
r80 68 88 0.326018
r81 67 83 0.652036
r82 67 68 15.6711
r83 66 69 0.655813
r84 65 88 0.326018
r85 65 66 4.58464
r86 48 79 1.82344
r87 43 57 1.16709
r88 43 73 2.16729
r89 38 69 1.82344
r90 35 48 1.16709
r91 30 38 1.16709
r92 25 57 0.0476429
r93 23 25 2.04225
r94 20 23 0.0685365
r95 18 23 0.5835
r96 18 19 2.8008
r97 15 19 0.652036
r98 8 20 3.8511
r99 6 35 0.185659
r100 4 15 3.8511
r101 2 30 0.185659
.ends

.subckt PM_G2_AOI21_N2_VDD 2 4 6 8 10 29 37 42 45 46 48 50 54 56 57 58 62 63 65
+ 67 68 74 Vss
c58 74 Vss 0.00462133f
c59 68 Vss 4.52364e-19
c60 65 Vss 0.00203839f
c61 63 Vss 0.00821501f
c62 62 Vss 8.61193e-19
c63 58 Vss 0.00179763f
c64 57 Vss 6.04409e-19
c65 56 Vss 0.00220637f
c66 54 Vss 0.00139836f
c67 51 Vss 0.00169975f
c68 50 Vss 0.0126653f
c69 48 Vss 0.00162243f
c70 46 Vss 0.00140335f
c71 45 Vss 0.00324454f
c72 42 Vss 0.00402078f
c73 37 Vss 0.00544429f
c74 33 Vss 0.0307649f
c75 29 Vss 1.05042e-19
c76 26 Vss 0.101606f
c77 22 Vss 0.035898f
c78 21 Vss 0.0712517f
c79 8 Vss 0.135377f
c80 6 Vss 0.136126f
c81 2 Vss 0.135008f
r82 64 68 0.551426
r83 64 65 4.58464
r84 63 68 0.551426
r85 62 67 0.326018
r86 62 63 15.5878
r87 58 68 0.0828784
r88 58 60 1.82344
r89 56 67 0.326018
r90 56 57 4.37625
r91 54 74 1.16709
r92 52 57 0.652036
r93 52 54 2.16729
r94 50 65 0.652036
r95 50 51 15.7128
r96 46 48 1.85991
r97 45 51 0.652036
r98 44 46 0.655813
r99 44 45 4.58464
r100 42 60 1.16709
r101 37 48 1.16709
r102 29 74 0.0476429
r103 27 33 0.494161
r104 27 29 1.45875
r105 26 30 0.652036
r106 26 29 1.45875
r107 23 33 0.128424
r108 21 33 0.494161
r109 21 22 2.8008
r110 18 22 0.652036
r111 10 42 0.185659
r112 8 30 3.8511
r113 6 23 3.8511
r114 4 37 0.185659
r115 2 18 3.8511
.ends

.subckt PM_G2_AOI21_N2_B 2 4 20 25 28 Vss
c17 28 Vss 0.00498247f
c18 25 Vss 6.10536e-19
c19 20 Vss 0.0915067f
c20 16 Vss 0.0598477f
c21 4 Vss 0.157143f
c22 2 Vss 0.372582f
r23 25 28 1.16709
r24 18 20 2.04225
r25 16 28 0.197068
r26 13 16 1.2837
r27 10 20 0.0685365
r28 8 18 0.0685365
r29 7 13 0.0685365
r30 4 10 4.3179
r31 2 8 9.9195
r32 2 7 3.8511
.ends

.subckt PM_G2_AOI21_N2_C 2 4 6 17 24 28 31 34 38 43 56 Vss
c46 56 Vss 0.00123749f
c47 43 Vss 0.0052622f
c48 38 Vss 0.00284502f
c49 34 Vss 0.00609886f
c50 28 Vss 0.0947914f
c51 24 Vss 0.0843207f
c52 17 Vss 3.53906e-19
c53 6 Vss 0.232307f
c54 4 Vss 0.201668f
c55 2 Vss 0.134559f
r56 52 56 0.652036
r57 38 56 5.16814
r58 34 43 1.16709
r59 34 52 10.4196
r60 31 34 0.145875
r61 26 28 2.04225
r62 24 43 0.0476429
r63 21 24 1.92555
r64 18 28 0.0685365
r65 17 38 1.16709
r66 13 26 0.0685365
r67 13 17 2.8008
r68 10 21 0.0685365
r69 6 18 7.1187
r70 4 17 4.3179
r71 2 10 3.8511
.ends

.subckt PM_G2_AOI21_N2_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00256251f
c33 27 Vss 0.00470045f
c34 23 Vss 0.00695334f
c35 8 Vss 0.00143442f
c36 6 Vss 0.00143442f
r37 33 35 7.002
r38 30 33 4.00114
r39 27 35 1.16709
r40 23 30 1.16709
r41 8 27 0.185659
r42 6 23 0.185659
r43 4 27 0.185659
r44 2 23 0.185659
.ends

.subckt PM_G2_AOI21_N2_A 2 4 10 11 13 14 15 20 24 29 32 Vss
c34 32 Vss 9.11501e-19
c35 29 Vss 4.23286e-19
c36 24 Vss 1.80739e-19
c37 20 Vss 0.136821f
c38 18 Vss 0.0247918f
c39 15 Vss 0.0322409f
c40 14 Vss 0.0730777f
c41 13 Vss 0.0312529f
c42 11 Vss 0.0324953f
c43 10 Vss 0.122088f
c44 2 Vss 0.238343f
r45 26 32 1.16709
r46 26 29 0.0729375
r47 24 32 0.262036
r48 20 32 0.238214
r49 18 24 0.326018
r50 18 20 0.64185
r51 15 24 2.50905
r52 14 24 0.326018
r53 14 24 0.1167
r54 13 15 0.652036
r55 12 13 1.22535
r56 10 12 0.652036
r57 10 11 3.09255
r58 7 11 0.652036
r59 4 20 3.7344
r60 2 7 7.4688
.ends

.subckt G2_AOI21_N2  VSS VDD B C Z A
*
* A	A
* Z	Z
* C	C
* B	B
* VDD	VDD
* VSS	VSS
XI14.X0 N_Z_XI14.X0_D N_VDD_XI14.X0_PGD N_A_XI14.X0_CG N_B_XI14.X0_PGS
+ N_VSS_XI14.X0_S TIGFET_HPNW8
XI12.X0 N_Z_XI12.X0_D N_VSS_XI12.X0_PGD N_B_XI12.X0_CG N_C_XI12.X0_PGS
+ N_VDD_XI12.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_VDD_XI15.X0_PGD N_C_XI15.X0_CG N_VDD_XI15.X0_PGS
+ N_VSS_XI15.X0_S TIGFET_HPNW8
XI13.X0 N_Z_XI13.X0_D N_VSS_XI13.X0_PGD N_A_XI13.X0_CG N_C_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW8
*
x_PM_G2_AOI21_N2_VSS N_VSS_XI14.X0_S N_VSS_XI12.X0_PGD N_VSS_XI15.X0_S
+ N_VSS_XI13.X0_PGD N_VSS_c_3_p N_VSS_c_35_p N_VSS_c_8_p N_VSS_c_2_p N_VSS_c_4_p
+ N_VSS_c_9_p N_VSS_c_5_p N_VSS_c_22_p N_VSS_c_10_p N_VSS_c_1_p N_VSS_c_6_p
+ N_VSS_c_7_p N_VSS_c_12_p N_VSS_c_15_p N_VSS_c_16_p VSS N_VSS_c_17_p Vss
+ PM_G2_AOI21_N2_VSS
x_PM_G2_AOI21_N2_VDD N_VDD_XI14.X0_PGD N_VDD_XI12.X0_S N_VDD_XI15.X0_PGD
+ N_VDD_XI15.X0_PGS N_VDD_XI13.X0_S N_VDD_c_80_p N_VDD_c_95_p N_VDD_c_96_p
+ N_VDD_c_79_p N_VDD_c_52_n N_VDD_c_53_n N_VDD_c_54_n N_VDD_c_74_p N_VDD_c_59_n
+ N_VDD_c_62_n N_VDD_c_63_n N_VDD_c_64_n N_VDD_c_65_n N_VDD_c_69_n VDD
+ N_VDD_c_72_n N_VDD_c_75_p Vss PM_G2_AOI21_N2_VDD
x_PM_G2_AOI21_N2_B N_B_XI14.X0_PGS N_B_XI12.X0_CG N_B_c_118_p B N_B_c_115_n Vss
+ PM_G2_AOI21_N2_B
x_PM_G2_AOI21_N2_C N_C_XI12.X0_PGS N_C_XI15.X0_CG N_C_XI13.X0_PGS N_C_c_139_n
+ N_C_c_142_n N_C_c_143_n C N_C_c_128_n N_C_c_131_n N_C_c_132_n N_C_c_136_n Vss
+ PM_G2_AOI21_N2_C
x_PM_G2_AOI21_N2_Z N_Z_XI14.X0_D N_Z_XI12.X0_D N_Z_XI15.X0_D N_Z_XI13.X0_D
+ N_Z_c_173_n N_Z_c_183_n N_Z_c_177_n Z Vss PM_G2_AOI21_N2_Z
x_PM_G2_AOI21_N2_A N_A_XI14.X0_CG N_A_XI13.X0_CG N_A_c_205_n N_A_c_217_n
+ N_A_c_218_n N_A_c_206_n N_A_c_219_n N_A_c_225_n N_A_c_207_n A N_A_c_210_n Vss
+ PM_G2_AOI21_N2_A
cc_1 N_VSS_c_1_p N_VDD_c_52_n 3.73937e-19
cc_2 N_VSS_c_2_p N_VDD_c_53_n 5.43852e-19
cc_3 N_VSS_c_3_p N_VDD_c_54_n 0.0012732f
cc_4 N_VSS_c_4_p N_VDD_c_54_n 0.00161703f
cc_5 N_VSS_c_5_p N_VDD_c_54_n 2.26455e-19
cc_6 N_VSS_c_6_p N_VDD_c_54_n 0.00447304f
cc_7 N_VSS_c_7_p N_VDD_c_54_n 0.00169823f
cc_8 N_VSS_c_8_p N_VDD_c_59_n 3.4118e-19
cc_9 N_VSS_c_9_p N_VDD_c_59_n 4.19648e-19
cc_10 N_VSS_c_10_p N_VDD_c_59_n 0.00353938f
cc_11 N_VSS_c_10_p N_VDD_c_62_n 0.00161744f
cc_12 N_VSS_c_12_p N_VDD_c_63_n 4.54377e-19
cc_13 N_VSS_c_10_p N_VDD_c_64_n 0.00106833f
cc_14 N_VSS_c_9_p N_VDD_c_65_n 0.00187494f
cc_15 N_VSS_c_15_p N_VDD_c_65_n 0.00340036f
cc_16 N_VSS_c_16_p N_VDD_c_65_n 0.00745699f
cc_17 N_VSS_c_17_p N_VDD_c_65_n 9.16632e-19
cc_18 N_VSS_c_4_p N_VDD_c_69_n 4.42007e-19
cc_19 N_VSS_c_5_p N_VDD_c_69_n 4.06699e-19
cc_20 N_VSS_c_16_p N_VDD_c_69_n 0.00303867f
cc_21 N_VSS_c_16_p N_VDD_c_72_n 0.00115015f
cc_22 N_VSS_c_22_p B 3.69138e-19
cc_23 N_VSS_c_10_p B 3.52052e-19
cc_24 N_VSS_XI12.X0_PGD N_C_XI12.X0_PGS 0.00151939f
cc_25 N_VSS_c_4_p N_C_c_128_n 8.90801e-19
cc_26 N_VSS_c_5_p N_C_c_128_n 3.44698e-19
cc_27 N_VSS_c_16_p N_C_c_128_n 0.00169235f
cc_28 N_VSS_c_16_p N_C_c_131_n 5.11302e-19
cc_29 N_VSS_XI12.X0_PGD N_C_c_132_n 3.23173e-19
cc_30 N_VSS_c_3_p N_C_c_132_n 0.00480946f
cc_31 N_VSS_c_4_p N_C_c_132_n 3.44698e-19
cc_32 N_VSS_c_5_p N_C_c_132_n 6.61756e-19
cc_33 N_VSS_c_10_p N_C_c_136_n 0.00251881f
cc_34 N_VSS_c_16_p N_C_c_136_n 3.90377e-19
cc_35 N_VSS_c_35_p N_Z_c_173_n 3.43419e-19
cc_36 N_VSS_c_8_p N_Z_c_173_n 3.43419e-19
cc_37 N_VSS_c_2_p N_Z_c_173_n 3.48267e-19
cc_38 N_VSS_c_9_p N_Z_c_173_n 3.48267e-19
cc_39 N_VSS_c_35_p N_Z_c_177_n 3.48267e-19
cc_40 N_VSS_c_8_p N_Z_c_177_n 3.48267e-19
cc_41 N_VSS_c_2_p N_Z_c_177_n 5.71987e-19
cc_42 N_VSS_c_9_p N_Z_c_177_n 5.71987e-19
cc_43 N_VSS_c_10_p N_Z_c_177_n 3.08274e-19
cc_44 N_VSS_c_16_p N_Z_c_177_n 7.49935e-19
cc_45 N_VSS_XI12.X0_PGD N_A_c_205_n 7.49544e-19
cc_46 N_VSS_XI13.X0_PGD N_A_c_206_n 0.00161855f
cc_47 N_VSS_c_5_p N_A_c_207_n 9.11194e-19
cc_48 N_VSS_c_4_p A 3.22909e-19
cc_49 N_VSS_c_5_p A 3.2351e-19
cc_50 N_VSS_c_4_p N_A_c_210_n 3.2351e-19
cc_51 N_VSS_c_5_p N_A_c_210_n 2.68747e-19
cc_52 N_VDD_XI14.X0_PGD N_B_XI14.X0_PGS 0.00174385f
cc_53 N_VDD_c_74_p B 6.29947e-19
cc_54 N_VDD_c_75_p B 3.48267e-19
cc_55 N_VDD_XI14.X0_PGD N_B_c_115_n 3.23173e-19
cc_56 N_VDD_c_74_p N_B_c_115_n 4.44903e-19
cc_57 N_VDD_c_75_p N_B_c_115_n 6.39485e-19
cc_58 N_VDD_c_79_p N_C_XI12.X0_PGS 2.86849e-19
cc_59 N_VDD_c_80_p N_C_c_139_n 9.37804e-19
cc_60 N_VDD_c_65_n N_C_c_139_n 5.88901e-19
cc_61 N_VDD_c_75_p N_C_c_139_n 2.68747e-19
cc_62 N_VDD_c_54_n N_C_c_142_n 3.8224e-19
cc_63 N_VDD_XI15.X0_PGS N_C_c_143_n 8.15793e-19
cc_64 N_VDD_c_65_n N_C_c_143_n 5.55843e-19
cc_65 N_VDD_c_79_p N_C_c_128_n 9.5543e-19
cc_66 N_VDD_c_53_n N_C_c_128_n 4.34676e-19
cc_67 N_VDD_c_54_n N_C_c_128_n 0.00198126f
cc_68 N_VDD_c_54_n N_C_c_131_n 6.31729e-19
cc_69 N_VDD_c_74_p N_C_c_131_n 4.21038e-19
cc_70 N_VDD_c_65_n N_C_c_131_n 4.49702e-19
cc_71 N_VDD_c_75_p N_C_c_131_n 3.2351e-19
cc_72 N_VDD_c_79_p N_C_c_132_n 3.63088e-19
cc_73 N_VDD_c_54_n N_C_c_132_n 2.64932e-19
cc_74 N_VDD_c_95_p N_Z_c_183_n 3.43419e-19
cc_75 N_VDD_c_96_p N_Z_c_183_n 3.43419e-19
cc_76 N_VDD_c_53_n N_Z_c_183_n 3.72424e-19
cc_77 N_VDD_c_54_n N_Z_c_183_n 3.4118e-19
cc_78 N_VDD_c_63_n N_Z_c_183_n 3.72199e-19
cc_79 N_VDD_c_95_p N_Z_c_177_n 3.48267e-19
cc_80 N_VDD_c_96_p N_Z_c_177_n 3.48267e-19
cc_81 N_VDD_c_53_n N_Z_c_177_n 5.09689e-19
cc_82 N_VDD_c_54_n N_Z_c_177_n 6.43655e-19
cc_83 N_VDD_c_63_n N_Z_c_177_n 7.72285e-19
cc_84 N_VDD_c_65_n N_Z_c_177_n 0.00139834f
cc_85 N_VDD_XI14.X0_PGD N_A_c_205_n 6.23873e-19
cc_86 N_VDD_XI15.X0_PGD N_A_c_206_n 3.69557e-19
cc_87 N_VDD_c_65_n A 4.8807e-19
cc_88 N_VDD_c_65_n N_A_c_210_n 3.66936e-19
cc_89 N_B_c_118_p N_C_XI12.X0_PGS 0.00196296f
cc_90 N_B_XI14.X0_PGS N_C_XI15.X0_CG 2.46172e-19
cc_91 N_B_c_118_p N_C_XI13.X0_PGS 4.66827e-19
cc_92 N_B_XI14.X0_PGS N_Z_c_177_n 2.61881e-19
cc_93 N_B_XI14.X0_PGS N_A_XI14.X0_CG 0.00881601f
cc_94 N_B_c_118_p N_A_c_217_n 0.00188162f
cc_95 N_B_XI14.X0_PGS N_A_c_218_n 6.07734e-19
cc_96 N_B_c_118_p N_A_c_219_n 0.00136534f
cc_97 N_B_c_118_p N_A_c_210_n 2.87722e-19
cc_98 N_C_c_139_n N_Z_c_177_n 9.83688e-19
cc_99 N_C_c_128_n N_Z_c_177_n 0.00274829f
cc_100 N_C_c_131_n N_Z_c_177_n 0.00329442f
cc_101 N_C_c_136_n N_Z_c_177_n 2.70867e-19
cc_102 N_C_XI15.X0_CG N_A_XI14.X0_CG 5.48933e-19
cc_103 N_C_c_139_n N_A_XI14.X0_CG 5.60239e-19
cc_104 N_C_XI13.X0_PGS N_A_c_205_n 8.10159e-19
cc_105 N_C_c_143_n N_A_c_205_n 0.00121323f
cc_106 N_C_XI13.X0_PGS N_A_c_225_n 4.5346e-19
cc_107 N_C_c_139_n N_A_c_207_n 9.47282e-19
cc_108 N_C_c_139_n A 4.56568e-19
cc_109 N_C_c_131_n A 6.34188e-19
cc_110 N_C_XI13.X0_PGS N_A_c_210_n 0.00570455f
cc_111 N_C_c_139_n N_A_c_210_n 6.1245e-19
cc_112 N_C_c_143_n N_A_c_210_n 0.00148932f
cc_113 N_C_c_131_n N_A_c_210_n 4.56568e-19
cc_114 N_Z_c_177_n N_A_XI14.X0_CG 5.52516e-19
cc_115 N_Z_c_173_n N_A_c_205_n 3.52706e-19
cc_116 N_Z_c_177_n N_A_c_205_n 3.09083e-19
cc_117 N_Z_c_183_n N_A_c_219_n 5.59623e-19
cc_118 N_Z_c_177_n A 0.00149422f
cc_119 N_Z_c_177_n N_A_c_210_n 9.63126e-19
*
.ends
*
*
.subckt AOI21_HPNW8 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 B0 Y A0) G2_AOI21_N2
.ends
*
* File: G2_BUF1_N2.pex.netlist
* Created: Wed Mar  2 15:38:39 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_BUF1_N2_VDD 2 4 7 11 28 30 32 44 48 52 54 56 57 61 65 67 71 75 78
+ 90 95 Vss
c59 95 Vss 0.0047576f
c60 90 Vss 0.00460635f
c61 80 Vss 9.22237e-19
c62 79 Vss 9.22237e-19
c63 75 Vss 0.00103298f
c64 71 Vss 9.84953e-19
c65 68 Vss 0.001766f
c66 67 Vss 0.0073616f
c67 65 Vss 0.00118372f
c68 61 Vss 0.00118372f
c69 57 Vss 0.00729501f
c70 56 Vss 0.0034296f
c71 54 Vss 0.00566164f
c72 52 Vss 0.0034296f
c73 51 Vss 0.001766f
c74 48 Vss 0.00382489f
c75 44 Vss 0.00532438f
c76 32 Vss 0.035607f
c77 31 Vss 0.102409f
c78 28 Vss 0.035607f
c79 27 Vss 0.102409f
c80 11 Vss 0.270897f
c81 7 Vss 0.270897f
r82 75 95 1.16709
r83 73 75 2.16729
r84 71 90 1.16709
r85 69 71 2.16729
r86 67 73 0.652036
r87 67 68 10.1279
r88 63 80 0.0828784
r89 63 65 1.82344
r90 59 79 0.0828784
r91 59 61 1.82344
r92 58 78 0.326018
r93 57 69 0.652036
r94 57 58 10.1279
r95 56 68 0.652036
r96 55 80 0.551426
r97 55 56 4.58464
r98 54 80 0.551426
r99 53 79 0.551426
r100 53 54 6.75193
r101 52 79 0.551426
r102 51 78 0.326018
r103 51 52 4.58464
r104 48 65 1.16709
r105 44 61 1.16709
r106 34 95 0.0476429
r107 32 34 1.45875
r108 31 38 0.652036
r109 31 34 1.45875
r110 30 90 0.0476429
r111 28 30 1.45875
r112 27 35 0.652036
r113 27 30 1.45875
r114 24 32 0.652036
r115 21 28 0.652036
r116 11 38 3.8511
r117 11 24 3.8511
r118 7 35 3.8511
r119 7 21 3.8511
r120 4 48 0.185659
r121 2 44 0.185659
.ends

.subckt PM_G2_BUF1_N2_VSS 3 7 10 12 27 28 30 31 32 45 49 52 57 62 67 72 77 97 98
+ 99 100 101 105 110 112 114 118 Vss
c56 116 Vss 6.78504e-19
c57 115 Vss 6.78504e-19
c58 114 Vss 0.00409661f
c59 112 Vss 0.00423582f
c60 110 Vss 0.0027381f
c61 105 Vss 0.0010217f
c62 101 Vss 8.62361e-19
c63 100 Vss 5.83649e-19
c64 99 Vss 0.00516968f
c65 98 Vss 5.83649e-19
c66 97 Vss 0.00631668f
c67 77 Vss 0.00400078f
c68 72 Vss 0.00410051f
c69 67 Vss 1.62518e-19
c70 62 Vss 7.10513e-22
c71 57 Vss 8.03422e-19
c72 52 Vss 9.77866e-19
c73 49 Vss 0.00537236f
c74 45 Vss 0.00387287f
c75 32 Vss 0.0350852f
c76 31 Vss 0.0994129f
c77 28 Vss 0.0350852f
c78 27 Vss 0.0994129f
c79 7 Vss 0.268864f
c80 3 Vss 0.268864f
r81 114 118 0.326018
r82 113 116 0.551426
r83 113 114 4.58464
r84 112 116 0.551426
r85 111 115 0.551426
r86 111 112 6.75193
r87 110 115 0.551426
r88 109 110 4.58464
r89 105 116 0.0828784
r90 101 115 0.0828784
r91 99 118 0.326018
r92 99 100 10.1279
r93 97 109 0.652036
r94 97 98 10.1279
r95 93 100 0.652036
r96 89 98 0.652036
r97 67 105 1.82344
r98 62 101 1.82344
r99 57 77 1.16709
r100 57 93 2.16729
r101 52 72 1.16709
r102 52 89 2.16729
r103 49 67 1.16709
r104 45 62 1.16709
r105 34 77 0.0476429
r106 32 34 1.45875
r107 31 38 0.652036
r108 31 34 1.45875
r109 30 72 0.0476429
r110 28 30 1.45875
r111 27 35 0.652036
r112 27 30 1.45875
r113 24 32 0.652036
r114 21 28 0.652036
r115 12 49 0.185659
r116 10 45 0.185659
r117 7 38 3.8511
r118 7 24 3.8511
r119 3 35 3.8511
r120 3 21 3.8511
.ends

.subckt PM_G2_BUF1_N2_A 2 4 12 22 28 Vss
c16 28 Vss 0.00294568f
c17 22 Vss 4.01518e-19
c18 12 Vss 0.200588f
c19 9 Vss 0.126125f
c20 7 Vss 0.0247918f
c21 4 Vss 0.139046f
r22 25 28 1.16709
r23 22 25 0.0416786
r24 15 28 0.0476429
r25 13 15 0.326018
r26 13 15 0.1167
r27 12 16 0.652036
r28 12 15 6.7686
r29 9 28 0.357321
r30 7 15 0.326018
r31 7 9 0.40845
r32 4 16 3.8511
r33 2 9 3.44265
.ends

.subckt PM_G2_BUF1_N2_Z 2 4 13 18 Vss
c14 18 Vss 4.84617e-19
c15 13 Vss 0.00522706f
c16 4 Vss 0.00176567f
r17 13 18 1.16709
r18 4 13 0.185659
r19 2 13 0.185659
.ends

.subckt PM_G2_BUF1_N2_NET17 2 4 6 8 18 33 36 41 50 58 Vss
c37 58 Vss 6.57973e-19
c38 50 Vss 0.00325633f
c39 41 Vss 0.00142824f
c40 36 Vss 0.00169654f
c41 33 Vss 0.00522706f
c42 22 Vss 0.0247918f
c43 19 Vss 0.0299669f
c44 18 Vss 0.169609f
c45 8 Vss 0.00176567f
c46 6 Vss 0.126125f
c47 2 Vss 0.138383f
r48 54 58 0.653045
r49 41 50 1.16709
r50 41 58 2.1395
r51 36 54 4.37625
r52 33 36 1.16709
r53 28 50 0.0476429
r54 26 50 0.357321
r55 22 28 0.326018
r56 22 26 0.40845
r57 19 28 6.7686
r58 18 28 0.326018
r59 18 28 0.1167
r60 15 19 0.652036
r61 8 33 0.185659
r62 6 26 3.44265
r63 4 33 0.185659
r64 2 15 3.8511
.ends

.subckt G2_BUF1_N2  VDD VSS A Z
*
* Z	Z
* A	A
* VSS	VSS
* VDD	VDD
XI10.X0 N_Z_XI10.X0_D N_VSS_XI10.X0_PGD N_NET17_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW8
XI7.X0 N_NET17_XI7.X0_D N_VSS_XI7.X0_PGD N_A_XI7.X0_CG N_VSS_XI7.X0_PGD
+ N_VDD_XI7.X0_S TIGFET_HPNW8
XI9.X0 N_Z_XI9.X0_D N_VDD_XI9.X0_PGD N_NET17_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW8
XI8.X0 N_NET17_XI8.X0_D N_VDD_XI8.X0_PGD N_A_XI8.X0_CG N_VDD_XI8.X0_PGD
+ N_VSS_XI8.X0_S TIGFET_HPNW8
*
x_PM_G2_BUF1_N2_VDD N_VDD_XI10.X0_S N_VDD_XI7.X0_S N_VDD_XI9.X0_PGD
+ N_VDD_XI8.X0_PGD N_VDD_c_4_p N_VDD_c_50_p N_VDD_c_8_p N_VDD_c_36_p
+ N_VDD_c_45_p N_VDD_c_6_p N_VDD_c_34_p N_VDD_c_3_p N_VDD_c_5_p N_VDD_c_38_p
+ N_VDD_c_46_p N_VDD_c_9_p N_VDD_c_13_p N_VDD_c_17_p VDD N_VDD_c_14_p
+ N_VDD_c_18_p Vss PM_G2_BUF1_N2_VDD
x_PM_G2_BUF1_N2_VSS N_VSS_XI10.X0_PGD N_VSS_XI7.X0_PGD N_VSS_XI9.X0_S
+ N_VSS_XI8.X0_S N_VSS_c_63_n N_VSS_c_65_n N_VSS_c_93_p N_VSS_c_67_n
+ N_VSS_c_69_n N_VSS_c_100_p N_VSS_c_106_p N_VSS_c_70_n N_VSS_c_74_n
+ N_VSS_c_101_p N_VSS_c_107_p N_VSS_c_78_n N_VSS_c_82_n N_VSS_c_85_n
+ N_VSS_c_86_n N_VSS_c_87_n N_VSS_c_88_n N_VSS_c_103_p N_VSS_c_110_p
+ N_VSS_c_89_n N_VSS_c_111_p N_VSS_c_90_n VSS Vss PM_G2_BUF1_N2_VSS
x_PM_G2_BUF1_N2_A N_A_XI7.X0_CG N_A_XI8.X0_CG N_A_c_116_n A N_A_c_119_n Vss
+ PM_G2_BUF1_N2_A
x_PM_G2_BUF1_N2_Z N_Z_XI10.X0_D N_Z_XI9.X0_D N_Z_c_132_n Z Vss PM_G2_BUF1_N2_Z
x_PM_G2_BUF1_N2_NET17 N_NET17_XI10.X0_CG N_NET17_XI7.X0_D N_NET17_XI9.X0_CG
+ N_NET17_XI8.X0_D N_NET17_c_147_n N_NET17_c_149_n N_NET17_c_151_n
+ N_NET17_c_154_n N_NET17_c_160_n N_NET17_c_163_n Vss PM_G2_BUF1_N2_NET17
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI10.X0_PGD 0.00201245f
cc_2 N_VDD_XI8.X0_PGD N_VSS_XI7.X0_PGD 0.00201245f
cc_3 N_VDD_c_3_p N_VSS_XI7.X0_PGD 3.05236e-19
cc_4 N_VDD_c_4_p N_VSS_c_63_n 0.00201245f
cc_5 N_VDD_c_5_p N_VSS_c_63_n 3.9313e-19
cc_6 N_VDD_c_6_p N_VSS_c_65_n 3.05236e-19
cc_7 N_VDD_c_5_p N_VSS_c_65_n 4.1253e-19
cc_8 N_VDD_c_8_p N_VSS_c_67_n 0.00201245f
cc_9 N_VDD_c_9_p N_VSS_c_67_n 3.9313e-19
cc_10 N_VDD_c_9_p N_VSS_c_69_n 4.1253e-19
cc_11 N_VDD_c_6_p N_VSS_c_70_n 8.67538e-19
cc_12 N_VDD_c_5_p N_VSS_c_70_n 0.00161703f
cc_13 N_VDD_c_13_p N_VSS_c_70_n 0.00106273f
cc_14 N_VDD_c_14_p N_VSS_c_70_n 3.48267e-19
cc_15 N_VDD_c_3_p N_VSS_c_74_n 8.67538e-19
cc_16 N_VDD_c_9_p N_VSS_c_74_n 0.00161703f
cc_17 N_VDD_c_17_p N_VSS_c_74_n 0.00110056f
cc_18 N_VDD_c_18_p N_VSS_c_74_n 3.48267e-19
cc_19 N_VDD_c_6_p N_VSS_c_78_n 3.66936e-19
cc_20 N_VDD_c_5_p N_VSS_c_78_n 2.26455e-19
cc_21 N_VDD_c_13_p N_VSS_c_78_n 3.99794e-19
cc_22 N_VDD_c_14_p N_VSS_c_78_n 6.489e-19
cc_23 N_VDD_c_3_p N_VSS_c_82_n 3.66936e-19
cc_24 N_VDD_c_9_p N_VSS_c_82_n 2.26455e-19
cc_25 N_VDD_c_18_p N_VSS_c_82_n 6.489e-19
cc_26 N_VDD_c_5_p N_VSS_c_85_n 0.00567457f
cc_27 N_VDD_c_5_p N_VSS_c_86_n 0.0017359f
cc_28 N_VDD_c_9_p N_VSS_c_87_n 0.00573644f
cc_29 N_VDD_c_9_p N_VSS_c_88_n 0.0017359f
cc_30 N_VDD_c_13_p N_VSS_c_89_n 3.85245e-19
cc_31 N_VDD_c_17_p N_VSS_c_90_n 3.85245e-19
cc_32 N_VDD_XI9.X0_PGD N_A_c_116_n 4.12647e-19
cc_33 N_VDD_XI8.X0_PGD N_A_c_116_n 4.07423e-19
cc_34 N_VDD_c_34_p A 9.3432e-19
cc_35 N_VDD_c_34_p N_A_c_119_n 5.18354e-19
cc_36 N_VDD_c_36_p N_Z_c_132_n 3.43419e-19
cc_37 N_VDD_c_5_p N_Z_c_132_n 3.4118e-19
cc_38 N_VDD_c_38_p N_Z_c_132_n 3.72199e-19
cc_39 N_VDD_c_36_p Z 3.48267e-19
cc_40 N_VDD_c_5_p Z 4.58391e-19
cc_41 N_VDD_c_38_p Z 7.4527e-19
cc_42 N_VDD_c_34_p N_NET17_XI10.X0_CG 2.86271e-19
cc_43 N_VDD_XI9.X0_PGD N_NET17_c_147_n 4.07423e-19
cc_44 N_VDD_XI8.X0_PGD N_NET17_c_147_n 4.12647e-19
cc_45 N_VDD_c_45_p N_NET17_c_149_n 3.43419e-19
cc_46 N_VDD_c_46_p N_NET17_c_149_n 3.72199e-19
cc_47 N_VDD_c_45_p N_NET17_c_151_n 3.48267e-19
cc_48 N_VDD_c_46_p N_NET17_c_151_n 8.0086e-19
cc_49 N_VDD_c_9_p N_NET17_c_151_n 4.34701e-19
cc_50 N_VDD_c_50_p N_NET17_c_154_n 3.02565e-19
cc_51 N_VDD_c_34_p N_NET17_c_154_n 2.74452e-19
cc_52 N_VDD_c_13_p N_NET17_c_154_n 4.44912e-19
cc_53 N_VDD_c_17_p N_NET17_c_154_n 2.83214e-19
cc_54 N_VDD_c_14_p N_NET17_c_154_n 3.49905e-19
cc_55 N_VDD_c_18_p N_NET17_c_154_n 4.45791e-19
cc_56 N_VDD_c_13_p N_NET17_c_160_n 3.43988e-19
cc_57 N_VDD_c_17_p N_NET17_c_160_n 2.24759e-19
cc_58 N_VDD_c_14_p N_NET17_c_160_n 2.68747e-19
cc_59 N_VDD_c_34_p N_NET17_c_163_n 4.34465e-19
cc_60 N_VSS_XI10.X0_PGD N_A_c_116_n 4.12647e-19
cc_61 N_VSS_XI7.X0_PGD N_A_c_116_n 4.04227e-19
cc_62 N_VSS_c_93_p A 2.23478e-19
cc_63 N_VSS_c_74_n A 3.28992e-19
cc_64 N_VSS_c_78_n A 2.26741e-19
cc_65 N_VSS_c_82_n A 6.58807e-19
cc_66 N_VSS_c_70_n N_A_c_119_n 2.11378e-19
cc_67 N_VSS_c_74_n N_A_c_119_n 3.2351e-19
cc_68 N_VSS_c_82_n N_A_c_119_n 2.68747e-19
cc_69 N_VSS_c_100_p N_Z_c_132_n 3.43419e-19
cc_70 N_VSS_c_101_p N_Z_c_132_n 3.48267e-19
cc_71 N_VSS_c_101_p Z 5.37696e-19
cc_72 N_VSS_c_103_p Z 2.7826e-19
cc_73 N_VSS_XI10.X0_PGD N_NET17_c_147_n 4.04227e-19
cc_74 N_VSS_XI7.X0_PGD N_NET17_c_147_n 4.12647e-19
cc_75 N_VSS_c_106_p N_NET17_c_149_n 3.43419e-19
cc_76 N_VSS_c_107_p N_NET17_c_149_n 3.48267e-19
cc_77 N_VSS_c_107_p N_NET17_c_151_n 4.8288e-19
cc_78 N_VSS_c_87_n N_NET17_c_151_n 4.84973e-19
cc_79 N_VSS_c_110_p N_NET17_c_151_n 5.49885e-19
cc_80 N_VSS_c_111_p N_NET17_c_151_n 0.00103514f
cc_81 N_VSS_c_85_n N_NET17_c_154_n 2.50699e-19
cc_82 N_VSS_c_111_p N_NET17_c_154_n 0.00119345f
cc_83 N_VSS_c_85_n N_NET17_c_163_n 8.43205e-19
cc_84 N_VSS_c_87_n N_NET17_c_163_n 4.88529e-19
cc_85 N_A_c_116_n N_NET17_c_147_n 0.0093393f
cc_86 N_A_c_116_n N_NET17_c_149_n 4.95639e-19
cc_87 A N_NET17_c_151_n 8.54729e-19
cc_88 N_Z_c_132_n N_NET17_c_147_n 4.95639e-19
cc_89 N_Z_c_132_n N_NET17_c_149_n 4.64289e-19
cc_90 Z N_NET17_c_149_n 2.11378e-19
cc_91 N_Z_c_132_n N_NET17_c_151_n 2.11378e-19
*
.ends
*
*
.subckt BUF1_HPNW8 A Y VDD VSS
xgate (VDD VSS A Y) G2_BUF1_N2
.ends
*
* File: G3_DFFQ1_N2.pex.netlist
* Created: Wed Apr  6 11:10:43 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_DFFQ1_N2_VSS 2 4 6 8 10 12 14 29 42 44 49 55 59 64 67 72 78 83 88
+ 93 102 111 116 125 126 127 128 132 137 142 148 154 156 161 163 165 166 167 Vss
c103 167 Vss 4.28045e-19
c104 166 Vss 3.75522e-19
c105 165 Vss 3.75522e-19
c106 164 Vss 6.15603e-19
c107 163 Vss 0.00495722f
c108 161 Vss 0.0016477f
c109 156 Vss 0.00136752f
c110 154 Vss 0.00253212f
c111 148 Vss 0.004602f
c112 142 Vss 0.00300844f
c113 132 Vss 0.0019674f
c114 128 Vss 6.73974e-19
c115 127 Vss 8.13835e-19
c116 126 Vss 0.00570183f
c117 125 Vss 0.00160501f
c118 116 Vss 0.00497548f
c119 111 Vss 0.00376876f
c120 102 Vss 0.00442938f
c121 93 Vss 2.73987e-19
c122 88 Vss 8.09754e-19
c123 83 Vss 7.28045e-19
c124 78 Vss 0.00155391f
c125 72 Vss 0.0108629f
c126 67 Vss 0.00135556f
c127 64 Vss 0.00650697f
c128 59 Vss 0.00498022f
c129 55 Vss 0.00373197f
c130 49 Vss 0.0568987f
c131 44 Vss 0.0568992f
c132 42 Vss 1.04992e-19
c133 29 Vss 0.035607f
c134 28 Vss 0.101294f
c135 14 Vss 0.134651f
c136 8 Vss 0.136772f
c137 6 Vss 0.133795f
c138 4 Vss 0.133902f
r139 162 167 0.551426
r140 162 163 15.5878
r141 161 167 0.551426
r142 160 161 4.62632
r143 156 167 0.0828784
r144 155 166 0.494161
r145 154 163 0.652036
r146 154 155 4.37625
r147 150 166 0.128424
r148 149 165 0.494161
r149 148 160 0.652036
r150 148 149 10.1279
r151 144 165 0.128424
r152 143 164 0.494161
r153 142 166 0.494161
r154 142 143 7.46046
r155 138 164 0.128424
r156 132 164 0.494161
r157 132 137 1.00029
r158 126 165 0.494161
r159 126 127 15.8795
r160 125 128 0.655813
r161 124 127 0.652036
r162 124 125 4.62632
r163 93 156 1.82344
r164 88 116 1.16709
r165 88 150 2.16729
r166 83 111 1.16709
r167 83 144 2.16729
r168 78 138 5.2515
r169 75 137 1.29204
r170 72 102 1.16709
r171 72 75 13.7539
r172 67 128 1.82344
r173 64 93 1.16709
r174 59 78 1.16709
r175 55 67 1.16709
r176 49 116 0.197068
r177 46 49 1.2837
r178 42 111 0.197068
r179 42 44 1.2837
r180 38 46 0.0685365
r181 35 44 0.0685365
r182 31 102 0.0476429
r183 29 31 1.45875
r184 28 32 0.652036
r185 28 31 1.45875
r186 25 29 0.652036
r187 14 38 3.8511
r188 12 64 0.185659
r189 10 59 0.185659
r190 8 35 3.8511
r191 6 32 3.8511
r192 4 25 3.8511
r193 2 55 0.185659
.ends

.subckt PM_G3_DFFQ1_N2_CK 2 4 6 8 18 21 25 37 40 Vss
c33 40 Vss 0.00476958f
c34 37 Vss 3.41336e-19
c35 33 Vss 0.0299314f
c36 25 Vss 0.166342f
c37 21 Vss 1.04992e-19
c38 18 Vss 0.18663f
c39 15 Vss 0.12596f
c40 13 Vss 0.0247918f
c41 6 Vss 0.550304f
c42 4 Vss 0.136627f
r43 37 40 1.16709
r44 26 33 0.494161
r45 25 27 0.652036
r46 25 26 4.84305
r47 22 33 0.128424
r48 21 40 0.0238214
r49 19 21 0.326018
r50 19 21 0.1167
r51 18 33 0.494161
r52 18 21 6.7686
r53 15 40 0.357321
r54 13 21 0.326018
r55 13 15 0.3501
r56 6 8 15.4044
r57 6 27 3.8511
r58 4 22 3.8511
r59 2 15 3.501
.ends

.subckt PM_G3_DFFQ1_N2_VDD 2 4 6 8 10 12 14 28 42 44 49 56 60 63 64 65 70 72 76
+ 78 79 82 84 86 91 93 95 96 98 99 100 102 104 113 118 Vss
c109 118 Vss 0.00535583f
c110 113 Vss 0.00546246f
c111 104 Vss 0.00475709f
c112 100 Vss 4.52364e-19
c113 99 Vss 2.39889e-19
c114 98 Vss 4.42806e-19
c115 96 Vss 0.00368915f
c116 95 Vss 5.05789e-19
c117 93 Vss 0.00304576f
c118 91 Vss 0.00856613f
c119 86 Vss 0.00179444f
c120 84 Vss 0.00304688f
c121 82 Vss 0.00102756f
c122 79 Vss 4.90412e-19
c123 78 Vss 0.00536329f
c124 76 Vss 6.6871e-19
c125 72 Vss 0.00341969f
c126 70 Vss 0.00232792f
c127 67 Vss 0.00182492f
c128 65 Vss 8.64465e-19
c129 64 Vss 0.00774944f
c130 63 Vss 0.00502551f
c131 60 Vss 0.00655192f
c132 56 Vss 0.00779243f
c133 49 Vss 0.0588939f
c134 44 Vss 0.0581359f
c135 42 Vss 1.01357e-19
c136 29 Vss 0.0372896f
c137 28 Vss 0.10099f
c138 12 Vss 0.13719f
c139 10 Vss 0.13484f
c140 8 Vss 0.00143442f
c141 4 Vss 0.136142f
c142 2 Vss 0.134971f
r143 95 104 1.16709
r144 95 96 0.470345
r145 93 102 0.326018
r146 92 100 0.551426
r147 92 93 4.58464
r148 91 100 0.551426
r149 90 91 15.6295
r150 86 100 0.0828784
r151 86 88 1.82344
r152 85 99 0.494161
r153 84 90 0.652036
r154 84 85 4.37625
r155 82 118 1.16709
r156 80 99 0.128424
r157 80 82 2.16729
r158 78 102 0.326018
r159 78 79 10.1279
r160 76 113 1.16709
r161 74 79 0.652036
r162 74 76 2.16729
r163 73 98 0.494161
r164 72 99 0.494161
r165 72 73 7.46046
r166 68 98 0.128424
r167 68 70 5.29318
r168 67 96 3.82922
r169 64 98 0.494161
r170 64 65 13.0037
r171 63 67 0.655813
r172 62 65 0.652036
r173 62 63 8.37739
r174 60 88 1.16709
r175 56 70 1.16709
r176 49 118 0.197068
r177 46 49 1.2837
r178 42 113 0.197068
r179 42 44 1.2837
r180 38 46 0.0685365
r181 35 44 0.0685365
r182 31 104 0.0476429
r183 29 31 1.45875
r184 28 32 0.652036
r185 28 31 1.45875
r186 25 29 0.652036
r187 14 60 0.185659
r188 12 38 3.8511
r189 10 35 3.8511
r190 8 56 0.185659
r191 6 56 0.185659
r192 4 25 3.8511
r193 2 32 3.8511
.ends

.subckt PM_G3_DFFQ1_N2_CKN 2 4 6 8 18 25 28 33 50 Vss
c38 51 Vss 0.00128326f
c39 50 Vss 0.00576518f
c40 33 Vss 7.37543e-19
c41 28 Vss 0.00177951f
c42 25 Vss 0.00542517f
c43 18 Vss 7.82969e-19
c44 6 Vss 0.475302f
c45 4 Vss 0.00143442f
r46 50 51 14.6709
r47 46 51 0.652036
r48 33 50 0.531835
r49 28 46 4.91807
r50 25 28 1.16709
r51 18 33 1.16709
r52 8 18 7.7022
r53 6 18 7.7022
r54 4 25 0.185659
r55 2 25 0.185659
.ends

.subckt PM_G3_DFFQ1_N2_D 2 4 11 12 22 25 28 Vss
c24 28 Vss 0.00170116f
c25 25 Vss 4.81931e-19
c26 12 Vss 0.21156f
c27 11 Vss 9.81474e-20
c28 7 Vss 0.0247918f
c29 4 Vss 0.137342f
c30 2 Vss 0.125849f
r31 25 28 1.16709
r32 22 25 0.0364688
r33 15 28 0.0476429
r34 13 15 0.326018
r35 13 15 0.1167
r36 12 16 0.652036
r37 12 15 6.7686
r38 11 28 0.357321
r39 7 15 0.326018
r40 7 11 0.40845
r41 4 16 3.8511
r42 2 11 3.44265
.ends

.subckt PM_G3_DFFQ1_N2_X 2 4 6 8 17 20 23 33 35 39 41 47 Vss
c47 47 Vss 0.00138877f
c48 41 Vss 5.3862e-19
c49 39 Vss 0.00123905f
c50 35 Vss 0.00217266f
c51 33 Vss 0.00551754f
c52 23 Vss 1.01432e-19
c53 20 Vss 0.21178f
c54 17 Vss 0.125802f
c55 15 Vss 0.0247918f
c56 8 Vss 0.137267f
c57 6 Vss 0.00143442f
r58 44 47 1.16709
r59 41 44 2.08393
r60 37 39 5.2515
r61 36 41 0.0685365
r62 35 37 0.652036
r63 35 36 1.70882
r64 33 39 1.16709
r65 23 47 0.0476429
r66 21 23 0.326018
r67 21 23 0.1167
r68 20 24 0.652036
r69 20 23 6.7686
r70 17 47 0.357321
r71 15 23 0.326018
r72 15 17 0.40845
r73 8 24 3.8511
r74 6 33 0.185659
r75 4 17 3.44265
r76 2 33 0.185659
.ends

.subckt PM_G3_DFFQ1_N2_Q 2 4 13 16 Vss
c12 16 Vss 3.81501e-19
c13 13 Vss 0.00450389f
c14 4 Vss 0.00143442f
r15 16 19 0.0416786
r16 13 19 1.16709
r17 4 13 0.185659
r18 2 13 0.185659
.ends

.subckt G3_DFFQ1_N2  VSS CK VDD D Q
*
* Q	Q
* D	D
* VDD	VDD
* CK	CK
* VSS	VSS
XI6.X0 N_CKN_XI6.X0_D N_VDD_XI6.X0_PGD N_CK_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW8
XI7.X0 N_CKN_XI7.X0_D N_VSS_XI7.X0_PGD N_CK_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW8
XI11.X0 N_X_XI11.X0_D N_VSS_XI11.X0_PGD N_D_XI11.X0_CG N_CK_XI11.X0_PGS
+ N_VDD_XI11.X0_S TIGFET_HPNW8
XI8.X0 N_Q_XI8.X0_D N_VDD_XI8.X0_PGD N_X_XI8.X0_CG N_CK_XI8.X0_PGS
+ N_VSS_XI8.X0_S TIGFET_HPNW8
XI10.X0 N_X_XI10.X0_D N_VDD_XI10.X0_PGD N_D_XI10.X0_CG N_CKN_XI10.X0_PGS
+ N_VSS_XI10.X0_S TIGFET_HPNW8
XI9.X0 N_Q_XI9.X0_D N_VSS_XI9.X0_PGD N_X_XI9.X0_CG N_CKN_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW8
*
x_PM_G3_DFFQ1_N2_VSS N_VSS_XI6.X0_S N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS
+ N_VSS_XI11.X0_PGD N_VSS_XI8.X0_S N_VSS_XI10.X0_S N_VSS_XI9.X0_PGD N_VSS_c_11_p
+ N_VSS_c_80_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_14_p N_VSS_c_101_p N_VSS_c_91_p
+ N_VSS_c_15_p N_VSS_c_3_p N_VSS_c_30_p N_VSS_c_21_p N_VSS_c_31_p N_VSS_c_41_p
+ N_VSS_c_53_p N_VSS_c_4_p N_VSS_c_34_p N_VSS_c_16_p N_VSS_c_7_p N_VSS_c_20_p
+ N_VSS_c_17_p N_VSS_c_77_p VSS N_VSS_c_35_p N_VSS_c_27_p N_VSS_c_36_p
+ N_VSS_c_43_p N_VSS_c_45_p N_VSS_c_46_p N_VSS_c_28_p N_VSS_c_37_p N_VSS_c_47_p
+ Vss PM_G3_DFFQ1_N2_VSS
x_PM_G3_DFFQ1_N2_CK N_CK_XI6.X0_CG N_CK_XI7.X0_CG N_CK_XI11.X0_PGS
+ N_CK_XI8.X0_PGS N_CK_c_108_n N_CK_c_125_p N_CK_c_109_n CK N_CK_c_115_p Vss
+ PM_G3_DFFQ1_N2_CK
x_PM_G3_DFFQ1_N2_VDD N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI7.X0_S
+ N_VDD_XI11.X0_S N_VDD_XI8.X0_PGD N_VDD_XI10.X0_PGD N_VDD_XI9.X0_S
+ N_VDD_c_140_n N_VDD_c_227_p N_VDD_c_141_n N_VDD_c_142_n N_VDD_c_214_p
+ N_VDD_c_240_p N_VDD_c_143_n N_VDD_c_147_n N_VDD_c_149_n N_VDD_c_150_n
+ N_VDD_c_152_n N_VDD_c_158_n N_VDD_c_161_n N_VDD_c_167_n N_VDD_c_168_n
+ N_VDD_c_170_n N_VDD_c_172_n N_VDD_c_173_n N_VDD_c_177_n N_VDD_c_181_n
+ N_VDD_c_183_n N_VDD_c_185_n N_VDD_c_186_n N_VDD_c_187_n VDD N_VDD_c_188_n
+ N_VDD_c_190_n N_VDD_c_193_n Vss PM_G3_DFFQ1_N2_VDD
x_PM_G3_DFFQ1_N2_CKN N_CKN_XI6.X0_D N_CKN_XI7.X0_D N_CKN_XI10.X0_PGS
+ N_CKN_XI9.X0_PGS N_CKN_c_261_n N_CKN_c_246_n N_CKN_c_248_n N_CKN_c_252_n
+ N_CKN_c_253_n Vss PM_G3_DFFQ1_N2_CKN
x_PM_G3_DFFQ1_N2_D N_D_XI11.X0_CG N_D_XI10.X0_CG N_D_c_284_n N_D_c_285_n D
+ N_D_c_286_n N_D_c_290_n Vss PM_G3_DFFQ1_N2_D
x_PM_G3_DFFQ1_N2_X N_X_XI11.X0_D N_X_XI8.X0_CG N_X_XI10.X0_D N_X_XI9.X0_CG
+ N_X_c_320_n N_X_c_308_n N_X_c_323_n N_X_c_309_n N_X_c_311_n N_X_c_312_n
+ N_X_c_316_n N_X_c_318_n Vss PM_G3_DFFQ1_N2_X
x_PM_G3_DFFQ1_N2_Q N_Q_XI8.X0_D N_Q_XI9.X0_D N_Q_c_355_n Q Vss PM_G3_DFFQ1_N2_Q
cc_1 N_VSS_XI7.X0_PGS N_CK_XI11.X0_PGS 0.00316278f
cc_2 N_VSS_XI11.X0_PGD N_CK_XI11.X0_PGS 0.00164185f
cc_3 N_VSS_c_3_p N_CK_XI11.X0_PGS 8.34822e-19
cc_4 N_VSS_c_4_p N_CK_XI11.X0_PGS 4.02129e-19
cc_5 N_VSS_XI7.X0_PGD N_CK_c_108_n 4.18808e-19
cc_6 N_VSS_XI7.X0_PGS N_CK_c_109_n 4.29708e-19
cc_7 N_VSS_c_7_p CK 5.33707e-19
cc_8 N_VSS_XI7.X0_PGD N_VDD_XI6.X0_PGD 0.00196344f
cc_9 N_VSS_XI9.X0_PGD N_VDD_XI8.X0_PGD 0.00221773f
cc_10 N_VSS_XI11.X0_PGD N_VDD_XI10.X0_PGD 0.00211593f
cc_11 N_VSS_c_11_p N_VDD_c_140_n 0.00196344f
cc_12 N_VSS_c_12_p N_VDD_c_141_n 0.00221773f
cc_13 N_VSS_c_13_p N_VDD_c_142_n 0.00211593f
cc_14 N_VSS_c_14_p N_VDD_c_143_n 9.5668e-19
cc_15 N_VSS_c_15_p N_VDD_c_143_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_143_n 0.00352032f
cc_17 N_VSS_c_17_p N_VDD_c_143_n 0.00185572f
cc_18 N_VSS_c_15_p N_VDD_c_147_n 4.50735e-19
cc_19 N_VSS_c_7_p N_VDD_c_147_n 0.00936712f
cc_20 N_VSS_c_20_p N_VDD_c_149_n 0.00105561f
cc_21 N_VSS_c_21_p N_VDD_c_150_n 0.00233232f
cc_22 N_VSS_c_4_p N_VDD_c_150_n 9.47758e-19
cc_23 N_VSS_c_13_p N_VDD_c_152_n 2.74851e-19
cc_24 N_VSS_c_21_p N_VDD_c_152_n 0.00161703f
cc_25 N_VSS_c_4_p N_VDD_c_152_n 2.24973e-19
cc_26 N_VSS_c_7_p N_VDD_c_152_n 0.00133545f
cc_27 N_VSS_c_27_p N_VDD_c_152_n 0.00408783f
cc_28 N_VSS_c_28_p N_VDD_c_152_n 7.74609e-19
cc_29 N_VSS_c_3_p N_VDD_c_158_n 0.00179097f
cc_30 N_VSS_c_30_p N_VDD_c_158_n 3.92901e-19
cc_31 N_VSS_c_31_p N_VDD_c_158_n 8.83788e-19
cc_32 N_VSS_c_12_p N_VDD_c_161_n 3.66315e-19
cc_33 N_VSS_c_31_p N_VDD_c_161_n 0.00141228f
cc_34 N_VSS_c_34_p N_VDD_c_161_n 0.00114511f
cc_35 N_VSS_c_35_p N_VDD_c_161_n 0.00409335f
cc_36 N_VSS_c_36_p N_VDD_c_161_n 0.00330569f
cc_37 N_VSS_c_37_p N_VDD_c_161_n 7.74609e-19
cc_38 N_VSS_c_35_p N_VDD_c_167_n 0.00144699f
cc_39 N_VSS_c_21_p N_VDD_c_168_n 9.29349e-19
cc_40 N_VSS_c_4_p N_VDD_c_168_n 3.79458e-19
cc_41 N_VSS_c_41_p N_VDD_c_170_n 4.50735e-19
cc_42 N_VSS_c_27_p N_VDD_c_170_n 0.00438429f
cc_43 N_VSS_c_43_p N_VDD_c_172_n 4.68065e-19
cc_44 N_VSS_c_41_p N_VDD_c_173_n 0.00187494f
cc_45 N_VSS_c_45_p N_VDD_c_173_n 0.00345634f
cc_46 N_VSS_c_46_p N_VDD_c_173_n 0.00778647f
cc_47 N_VSS_c_47_p N_VDD_c_173_n 9.16632e-19
cc_48 N_VSS_c_31_p N_VDD_c_177_n 4.35319e-19
cc_49 N_VSS_c_34_p N_VDD_c_177_n 3.66936e-19
cc_50 N_VSS_c_36_p N_VDD_c_177_n 0.00106857f
cc_51 N_VSS_c_46_p N_VDD_c_177_n 0.00335989f
cc_52 N_VSS_c_3_p N_VDD_c_181_n 6.19689e-19
cc_53 N_VSS_c_53_p N_VDD_c_181_n 3.8721e-19
cc_54 N_VSS_c_15_p N_VDD_c_183_n 0.00222015f
cc_55 N_VSS_c_7_p N_VDD_c_183_n 2.66524e-19
cc_56 N_VSS_c_7_p N_VDD_c_185_n 0.00118128f
cc_57 N_VSS_c_27_p N_VDD_c_186_n 0.0010448f
cc_58 N_VSS_c_46_p N_VDD_c_187_n 0.00116512f
cc_59 N_VSS_c_3_p N_VDD_c_188_n 3.86162e-19
cc_60 N_VSS_c_53_p N_VDD_c_188_n 6.0892e-19
cc_61 N_VSS_c_3_p N_VDD_c_190_n 5.2607e-19
cc_62 N_VSS_c_31_p N_VDD_c_190_n 3.48267e-19
cc_63 N_VSS_c_34_p N_VDD_c_190_n 6.489e-19
cc_64 N_VSS_c_21_p N_VDD_c_193_n 3.48267e-19
cc_65 N_VSS_c_4_p N_VDD_c_193_n 6.20986e-19
cc_66 N_VSS_c_14_p N_CKN_c_246_n 3.43419e-19
cc_67 N_VSS_c_15_p N_CKN_c_246_n 3.48267e-19
cc_68 N_VSS_c_15_p N_CKN_c_248_n 0.00109746f
cc_69 N_VSS_c_3_p N_CKN_c_248_n 6.97825e-19
cc_70 N_VSS_c_7_p N_CKN_c_248_n 4.81255e-19
cc_71 N_VSS_c_46_p N_CKN_c_248_n 2.6973e-19
cc_72 N_VSS_c_46_p N_CKN_c_252_n 0.00111539f
cc_73 N_VSS_c_3_p N_CKN_c_253_n 0.00225294f
cc_74 N_VSS_c_30_p N_CKN_c_253_n 7.04847e-19
cc_75 N_VSS_c_31_p N_CKN_c_253_n 6.45464e-19
cc_76 N_VSS_c_7_p N_CKN_c_253_n 0.00132819f
cc_77 N_VSS_c_77_p N_CKN_c_253_n 7.24142e-19
cc_78 N_VSS_c_35_p N_CKN_c_253_n 7.58219e-19
cc_79 N_VSS_c_27_p N_CKN_c_253_n 9.23091e-19
cc_80 N_VSS_c_80_p N_D_c_284_n 9.24646e-19
cc_81 N_VSS_XI11.X0_PGD N_D_c_285_n 3.94389e-19
cc_82 N_VSS_c_3_p N_D_c_286_n 6.13924e-19
cc_83 N_VSS_c_21_p N_D_c_286_n 2.96367e-19
cc_84 N_VSS_c_53_p N_D_c_286_n 3.48267e-19
cc_85 N_VSS_c_4_p N_D_c_286_n 3.20302e-19
cc_86 N_VSS_c_3_p N_D_c_290_n 3.48267e-19
cc_87 N_VSS_c_21_p N_D_c_290_n 3.20302e-19
cc_88 N_VSS_c_53_p N_D_c_290_n 6.88619e-19
cc_89 N_VSS_c_4_p N_D_c_290_n 2.62417e-19
cc_90 N_VSS_XI9.X0_PGD N_X_c_308_n 4.04227e-19
cc_91 N_VSS_c_91_p N_X_c_309_n 3.43419e-19
cc_92 N_VSS_c_41_p N_X_c_309_n 3.48267e-19
cc_93 N_VSS_c_35_p N_X_c_311_n 2.44303e-19
cc_94 N_VSS_c_91_p N_X_c_312_n 3.48267e-19
cc_95 N_VSS_c_3_p N_X_c_312_n 4.71026e-19
cc_96 N_VSS_c_41_p N_X_c_312_n 5.71987e-19
cc_97 N_VSS_c_46_p N_X_c_312_n 2.97611e-19
cc_98 N_VSS_c_3_p N_X_c_316_n 0.00157847f
cc_99 N_VSS_c_46_p N_X_c_316_n 2.88807e-19
cc_100 N_VSS_c_3_p N_X_c_318_n 3.48267e-19
cc_101 N_VSS_c_101_p N_Q_c_355_n 3.43419e-19
cc_102 N_VSS_c_30_p N_Q_c_355_n 3.48267e-19
cc_103 N_VSS_c_30_p Q 5.37696e-19
cc_104 N_CK_c_108_n N_VDD_XI6.X0_PGD 4.18808e-19
cc_105 N_CK_XI11.X0_PGS N_VDD_XI10.X0_PGD 2.44781e-19
cc_106 N_CK_c_109_n N_VDD_c_142_n 2.44781e-19
cc_107 CK N_VDD_c_143_n 5.04211e-19
cc_108 N_CK_c_115_p N_VDD_c_143_n 5.30123e-19
cc_109 N_CK_c_108_n N_VDD_c_147_n 0.0015171f
cc_110 CK N_VDD_c_147_n 0.00141439f
cc_111 N_CK_c_115_p N_VDD_c_147_n 0.00120239f
cc_112 N_CK_XI11.X0_PGS N_VDD_c_150_n 2.48209e-19
cc_113 N_CK_c_109_n N_VDD_c_150_n 5.56076e-19
cc_114 CK N_VDD_c_150_n 3.85155e-19
cc_115 N_CK_c_115_p N_VDD_c_150_n 2.72301e-19
cc_116 CK N_VDD_c_181_n 4.2144e-19
cc_117 N_CK_c_115_p N_VDD_c_181_n 3.27641e-19
cc_118 N_CK_c_125_p N_VDD_c_188_n 9.40274e-19
cc_119 CK N_VDD_c_188_n 3.20302e-19
cc_120 N_CK_c_115_p N_VDD_c_188_n 2.62417e-19
cc_121 N_CK_XI11.X0_PGS N_CKN_XI10.X0_PGS 4.11563e-19
cc_122 N_CK_XI11.X0_PGS N_CKN_c_261_n 2.73384e-19
cc_123 N_CK_c_108_n N_CKN_c_246_n 6.55689e-19
cc_124 N_CK_XI11.X0_PGS N_D_XI11.X0_CG 4.28946e-19
cc_125 N_CK_XI11.X0_PGS N_D_XI10.X0_CG 2.59344e-19
cc_126 N_CK_XI11.X0_PGS N_D_c_290_n 0.00300565f
cc_127 N_CK_XI11.X0_PGS N_X_XI9.X0_CG 2.61247e-19
cc_128 N_CK_XI11.X0_PGS N_X_c_320_n 4.55333e-19
cc_129 N_CK_XI11.X0_PGS N_X_c_318_n 0.00630896f
cc_130 N_VDD_c_173_n N_CKN_XI10.X0_PGS 7.25969e-19
cc_131 N_VDD_c_173_n N_CKN_c_261_n 8.21431e-19
cc_132 N_VDD_c_214_p N_CKN_c_246_n 3.43419e-19
cc_133 N_VDD_c_214_p N_CKN_c_248_n 3.48267e-19
cc_134 N_VDD_c_143_n N_CKN_c_248_n 3.84058e-19
cc_135 N_VDD_c_147_n N_CKN_c_248_n 4.28606e-19
cc_136 N_VDD_c_150_n N_CKN_c_248_n 5.37696e-19
cc_137 N_VDD_c_181_n N_CKN_c_248_n 6.42405e-19
cc_138 N_VDD_c_173_n N_CKN_c_252_n 7.71262e-19
cc_139 N_VDD_c_147_n N_CKN_c_253_n 3.98085e-19
cc_140 N_VDD_c_152_n N_CKN_c_253_n 2.80228e-19
cc_141 N_VDD_c_161_n N_CKN_c_253_n 4.0976e-19
cc_142 N_VDD_c_168_n N_CKN_c_253_n 2.45963e-19
cc_143 N_VDD_XI10.X0_PGD N_D_c_285_n 4.07433e-19
cc_144 N_VDD_XI8.X0_PGD N_X_c_308_n 3.96342e-19
cc_145 N_VDD_c_227_p N_X_c_323_n 8.75838e-19
cc_146 N_VDD_c_214_p N_X_c_309_n 3.43419e-19
cc_147 N_VDD_c_150_n N_X_c_309_n 3.48267e-19
cc_148 N_VDD_c_152_n N_X_c_309_n 3.37713e-19
cc_149 N_VDD_c_214_p N_X_c_312_n 3.48267e-19
cc_150 N_VDD_c_150_n N_X_c_312_n 6.94315e-19
cc_151 N_VDD_c_152_n N_X_c_312_n 4.72817e-19
cc_152 N_VDD_c_173_n N_X_c_312_n 0.00111552f
cc_153 N_VDD_c_158_n N_X_c_316_n 4.35824e-19
cc_154 N_VDD_c_173_n N_X_c_316_n 2.02855e-19
cc_155 N_VDD_c_190_n N_X_c_316_n 3.40502e-19
cc_156 N_VDD_c_158_n N_X_c_318_n 3.43988e-19
cc_157 N_VDD_c_190_n N_X_c_318_n 2.68747e-19
cc_158 N_VDD_c_240_p N_Q_c_355_n 3.43419e-19
cc_159 N_VDD_c_161_n N_Q_c_355_n 3.4118e-19
cc_160 N_VDD_c_172_n N_Q_c_355_n 3.72199e-19
cc_161 N_VDD_c_240_p Q 3.48267e-19
cc_162 N_VDD_c_161_n Q 4.58391e-19
cc_163 N_VDD_c_172_n Q 7.06537e-19
cc_164 N_CKN_XI10.X0_PGS N_D_XI10.X0_CG 0.00419505f
cc_165 N_CKN_XI10.X0_PGS N_X_c_308_n 0.00425073f
cc_166 N_CKN_c_261_n N_X_c_311_n 5.71169e-19
cc_167 N_CKN_c_253_n N_X_c_311_n 0.00127072f
cc_168 N_CKN_c_248_n N_X_c_312_n 4.96487e-19
cc_169 N_CKN_c_252_n N_X_c_312_n 8.08281e-19
cc_170 N_CKN_c_253_n N_X_c_312_n 6.84099e-19
cc_171 N_CKN_c_253_n N_X_c_316_n 8.25313e-19
cc_172 N_D_c_285_n N_X_c_308_n 0.00474388f
cc_173 N_D_c_285_n N_X_c_309_n 6.8653e-19
cc_174 N_D_c_285_n N_X_c_312_n 3.40033e-19
cc_175 N_D_c_286_n N_X_c_312_n 0.00151909f
cc_176 N_D_c_290_n N_X_c_312_n 0.00104518f
cc_177 N_D_c_286_n N_X_c_316_n 0.00146206f
cc_178 N_D_c_290_n N_X_c_316_n 0.00103457f
cc_179 N_D_c_286_n N_X_c_318_n 4.56568e-19
cc_180 N_D_c_290_n N_X_c_318_n 0.00373359f
cc_181 N_X_c_308_n N_Q_c_355_n 6.8653e-19
cc_182 N_X_c_311_n N_Q_c_355_n 4.47287e-19
cc_183 N_X_c_311_n Q 6.7453e-19
*
.ends
*
*
.subckt DFFQ1_HPNW8 CK D Q VDD VSS
xgate (VSS CK VDD D Q) G3_DFFQ1_N2
.ends
*
* File: G1_INV1_N2.pex.netlist
* Created: Fri Feb 25 16:24:20 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G1_INV1_N2_VDD 2 5 15 23 28 30 34 37 43 Vss
c22 43 Vss 0.00440656f
c23 34 Vss 7.98732e-19
c24 30 Vss 0.00489873f
c25 28 Vss 0.00252866f
c26 26 Vss 0.00167653f
c27 23 Vss 0.00387287f
c28 15 Vss 0.035607f
c29 14 Vss 0.102409f
c30 5 Vss 0.271444f
r31 34 43 1.16709
r32 32 34 2.41736
r33 31 37 0.326018
r34 30 32 0.652036
r35 30 31 7.46046
r36 26 37 0.326018
r37 26 28 5.50157
r38 23 28 1.16709
r39 17 43 0.0476429
r40 15 17 1.45875
r41 14 18 0.652036
r42 14 17 1.45875
r43 11 15 0.652036
r44 5 18 3.8511
r45 5 11 3.8511
r46 2 23 0.185659
.ends

.subckt PM_G1_INV1_N2_A 2 4 12 22 25 28 Vss
c7 28 Vss 0.00718398f
c8 12 Vss 0.22585f
c9 9 Vss 0.126125f
c10 7 Vss 0.0247918f
c11 4 Vss 0.139046f
r12 22 28 1.16709
r13 22 25 0.0416786
r14 15 28 0.0476429
r15 13 15 0.326018
r16 13 15 0.1167
r17 12 16 0.652036
r18 12 15 6.7686
r19 9 28 0.357321
r20 7 15 0.326018
r21 7 9 0.40845
r22 4 16 3.8511
r23 2 9 3.44265
.ends

.subckt PM_G1_INV1_N2_VSS 3 6 14 24 27 32 37 49 50 56 Vss
c24 51 Vss 0.0012655f
c25 50 Vss 6.56963e-19
c26 49 Vss 0.00353949f
c27 37 Vss 0.00375421f
c28 32 Vss 0.00198022f
c29 27 Vss 2.9624e-19
c30 24 Vss 0.00537236f
c31 15 Vss 0.0358979f
c32 14 Vss 0.0994171f
c33 3 Vss 0.270557f
r34 51 56 0.326018
r35 49 56 0.326018
r36 49 50 7.46046
r37 45 50 0.652036
r38 32 51 5.50157
r39 27 37 1.16709
r40 27 45 2.41736
r41 24 32 1.16709
r42 17 37 0.0476429
r43 15 17 1.45875
r44 14 18 0.652036
r45 14 17 1.45875
r46 11 15 0.652036
r47 6 24 0.185659
r48 3 18 3.8511
r49 3 11 3.8511
.ends

.subckt PM_G1_INV1_N2_Z 2 4 13 16 Vss
c11 13 Vss 0.00523231f
c12 4 Vss 0.00143442f
r13 16 19 0.0416786
r14 13 19 1.16709
r15 4 13 0.185659
r16 2 13 0.185659
.ends

.subckt G1_INV1_N2  VDD A VSS Z
*
* Z	Z
* VSS	VSS
* A	A
* VDD	VDD
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_A_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VDD_XI4.X0_PGD N_A_XI4.X0_CG N_VDD_XI4.X0_PGD
+ N_VSS_XI4.X0_S TIGFET_HPNW8
*
x_PM_G1_INV1_N2_VDD N_VDD_XI6.X0_S N_VDD_XI4.X0_PGD N_VDD_c_4_p N_VDD_c_17_p
+ N_VDD_c_3_p N_VDD_c_5_p N_VDD_c_8_p VDD N_VDD_c_9_p Vss PM_G1_INV1_N2_VDD
x_PM_G1_INV1_N2_A N_A_XI6.X0_CG N_A_XI4.X0_CG N_A_c_23_n N_A_c_25_p A N_A_c_26_p
+ Vss PM_G1_INV1_N2_A
x_PM_G1_INV1_N2_VSS N_VSS_XI6.X0_PGD N_VSS_XI4.X0_S N_VSS_c_32_n N_VSS_c_50_p
+ N_VSS_c_34_n N_VSS_c_38_n N_VSS_c_40_n N_VSS_c_43_n N_VSS_c_44_n VSS Vss
+ PM_G1_INV1_N2_VSS
x_PM_G1_INV1_N2_Z N_Z_XI6.X0_D N_Z_XI4.X0_D N_Z_c_54_n Z Vss PM_G1_INV1_N2_Z
cc_1 N_VDD_XI4.X0_PGD N_A_c_23_n 4.28964e-19
cc_2 N_VDD_XI4.X0_PGD N_VSS_XI6.X0_PGD 0.0020004f
cc_3 N_VDD_c_3_p N_VSS_XI6.X0_PGD 4.31044e-19
cc_4 N_VDD_c_4_p N_VSS_c_32_n 0.0020004f
cc_5 N_VDD_c_5_p N_VSS_c_32_n 5.13652e-19
cc_6 N_VDD_c_3_p N_VSS_c_34_n 0.00287439f
cc_7 N_VDD_c_5_p N_VSS_c_34_n 0.00141709f
cc_8 N_VDD_c_8_p N_VSS_c_34_n 8.61874e-19
cc_9 N_VDD_c_9_p N_VSS_c_34_n 3.48267e-19
cc_10 N_VDD_c_3_p N_VSS_c_38_n 4.56935e-19
cc_11 N_VDD_c_8_p N_VSS_c_38_n 0.00104259f
cc_12 N_VDD_c_3_p N_VSS_c_40_n 9.55109e-19
cc_13 N_VDD_c_5_p N_VSS_c_40_n 0.00103739f
cc_14 N_VDD_c_9_p N_VSS_c_40_n 6.46219e-19
cc_15 N_VDD_c_5_p N_VSS_c_43_n 0.00582834f
cc_16 N_VDD_c_5_p N_VSS_c_44_n 0.00172765f
cc_17 N_VDD_c_17_p N_Z_c_54_n 3.43419e-19
cc_18 N_VDD_c_3_p N_Z_c_54_n 3.48267e-19
cc_19 N_VDD_c_5_p N_Z_c_54_n 3.21105e-19
cc_20 N_VDD_c_17_p Z 3.48267e-19
cc_21 N_VDD_c_3_p Z 7.09569e-19
cc_22 N_VDD_c_5_p Z 4.30066e-19
cc_23 N_A_c_23_n N_VSS_XI6.X0_PGD 4.2599e-19
cc_24 N_A_c_25_p N_VSS_c_34_n 6.08006e-19
cc_25 N_A_c_26_p N_VSS_c_34_n 3.34201e-19
cc_26 N_A_c_25_p N_VSS_c_40_n 3.49905e-19
cc_27 N_A_c_26_p N_VSS_c_40_n 2.68747e-19
cc_28 N_A_c_23_n N_Z_c_54_n 6.55689e-19
cc_29 N_VSS_c_50_p N_Z_c_54_n 3.43419e-19
cc_30 N_VSS_c_38_n N_Z_c_54_n 3.48267e-19
cc_31 N_VSS_c_38_n Z 8.23589e-19
cc_32 N_VSS_c_43_n Z 2.41335e-19
*
.ends
*
*
.subckt INV1_HPNW8 A Y VDD VSS
xgate (VDD A VSS Y) G1_INV1_N2
.ends
*
* File: G3_LATQ1_N2.pex.netlist
* Created: Tue Apr  5 11:38:39 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_LATQ1_N2_VDD 2 4 6 8 10 12 14 16 31 42 44 48 58 63 66 68 69 70 71
+ 72 75 77 81 85 90 92 98 103 Vss
c89 103 Vss 0.00490183f
c90 98 Vss 0.00460926f
c91 90 Vss 2.39889e-19
c92 85 Vss 0.00243594f
c93 83 Vss 0.0016991f
c94 81 Vss 9.06638e-19
c95 77 Vss 0.0042879f
c96 75 Vss 7.26394e-19
c97 72 Vss 8.65068e-19
c98 71 Vss 0.0022063f
c99 70 Vss 8.64091e-19
c100 69 Vss 0.00567616f
c101 68 Vss 0.00905486f
c102 66 Vss 0.00502493f
c103 63 Vss 0.00660615f
c104 58 Vss 0.00394659f
c105 53 Vss 0.0307649f
c106 48 Vss 0.231494f
c107 44 Vss 7.7692e-20
c108 42 Vss 0.0357051f
c109 41 Vss 0.0656875f
c110 32 Vss 0.035919f
c111 31 Vss 0.101295f
c112 16 Vss 0.00143442f
c113 14 Vss 0.137165f
c114 10 Vss 0.136745f
c115 8 Vss 0.135164f
c116 6 Vss 0.13553f
c117 4 Vss 0.135175f
r118 83 92 0.326018
r119 83 85 5.2515
r120 81 103 1.16709
r121 79 81 2.16729
r122 78 90 0.494161
r123 77 92 0.326018
r124 77 78 7.46046
r125 75 98 1.16709
r126 73 90 0.128424
r127 73 75 2.16729
r128 71 90 0.494161
r129 71 72 4.37625
r130 69 79 0.652036
r131 69 70 10.1279
r132 68 72 0.652036
r133 67 68 15.5461
r134 66 89 2.334
r135 66 67 0.14525
r136 65 70 0.652036
r137 65 66 4.62632
r138 63 85 1.16709
r139 58 89 1.16709
r140 49 53 0.494161
r141 48 50 0.652036
r142 48 49 6.8853
r143 45 53 0.128424
r144 44 103 0.0476429
r145 42 44 1.45875
r146 41 53 0.494161
r147 41 44 1.45875
r148 38 42 0.652036
r149 34 98 0.0476429
r150 32 34 1.45875
r151 31 35 0.652036
r152 31 34 1.45875
r153 28 32 0.652036
r154 16 63 0.185659
r155 14 50 3.8511
r156 12 63 0.185659
r157 10 45 3.8511
r158 8 38 3.8511
r159 6 28 3.8511
r160 4 35 3.8511
r161 2 58 0.185659
.ends

.subckt PM_G3_LATQ1_N2_VSS 2 4 6 8 10 12 14 16 31 32 34 42 48 58 63 66 71 76 81
+ 90 95 104 106 107 108 113 114 119 129 130 132 Vss
c81 130 Vss 3.75522e-19
c82 129 Vss 4.28045e-19
c83 125 Vss 0.00128107f
c84 119 Vss 0.00326562f
c85 114 Vss 8.21919e-19
c86 113 Vss 0.00415461f
c87 108 Vss 8.27105e-19
c88 107 Vss 0.00171853f
c89 106 Vss 0.00164009f
c90 104 Vss 0.00508678f
c91 95 Vss 0.00436437f
c92 90 Vss 0.00392783f
c93 81 Vss 0.0023337f
c94 76 Vss 5.9672e-19
c95 71 Vss 4.65089e-19
c96 66 Vss 0.00142325f
c97 63 Vss 0.00655541f
c98 58 Vss 0.00751018f
c99 53 Vss 0.0307649f
c100 48 Vss 0.231624f
c101 42 Vss 0.0348714f
c102 41 Vss 0.0648006f
c103 34 Vss 1.05421e-19
c104 32 Vss 0.0350852f
c105 31 Vss 0.0994129f
c106 16 Vss 0.137353f
c107 14 Vss 0.00143442f
c108 12 Vss 0.137077f
c109 10 Vss 0.135163f
c110 4 Vss 0.135531f
c111 2 Vss 0.135176f
r112 125 132 0.326018
r113 120 130 0.494161
r114 119 132 0.326018
r115 119 120 7.46046
r116 115 130 0.128424
r117 113 121 0.652036
r118 113 114 10.1279
r119 109 129 0.0828784
r120 107 130 0.494161
r121 107 108 4.37625
r122 106 114 0.652036
r123 105 129 0.551426
r124 105 106 4.58464
r125 104 129 0.551426
r126 103 108 0.652036
r127 103 104 15.5878
r128 81 125 5.2515
r129 76 95 1.16709
r130 76 121 2.16729
r131 71 90 1.16709
r132 71 115 2.16729
r133 66 109 1.82344
r134 63 81 1.16709
r135 58 66 1.16709
r136 49 53 0.494161
r137 48 50 0.652036
r138 48 49 6.8853
r139 45 53 0.128424
r140 44 95 0.0476429
r141 42 44 1.45875
r142 41 53 0.494161
r143 41 44 1.45875
r144 38 42 0.652036
r145 34 90 0.0476429
r146 32 34 1.45875
r147 31 35 0.652036
r148 31 34 1.45875
r149 28 32 0.652036
r150 16 50 3.8511
r151 14 63 0.185659
r152 12 45 3.8511
r153 10 38 3.8511
r154 8 63 0.185659
r155 6 58 0.185659
r156 4 28 3.8511
r157 2 35 3.8511
.ends

.subckt PM_G3_LATQ1_N2_G 2 4 6 14 15 22 31 37 Vss
c26 37 Vss 0.00234039f
c27 31 Vss 4.77975e-19
c28 29 Vss 0.0295006f
c29 22 Vss 0.152742f
c30 15 Vss 0.17649f
c31 14 Vss 2.16373e-19
c32 10 Vss 0.0247918f
c33 6 Vss 0.137829f
c34 4 Vss 0.138596f
c35 2 Vss 0.125945f
r36 34 37 1.16709
r37 31 34 0.0833571
r38 23 29 0.494161
r39 22 24 0.652036
r40 22 23 4.84305
r41 19 29 0.128424
r42 18 37 0.0476429
r43 16 18 0.326018
r44 16 18 0.1167
r45 15 29 0.494161
r46 15 18 6.7686
r47 14 37 0.357321
r48 10 18 0.326018
r49 10 14 0.40845
r50 6 24 3.8511
r51 4 19 3.8511
r52 2 14 3.44265
.ends

.subckt PM_G3_LATQ1_N2_QN 2 4 6 8 20 23 33 37 40 45 48 53 69 Vss
c46 69 Vss 4.0109e-19
c47 53 Vss 0.0021144f
c48 48 Vss 0.00823447f
c49 45 Vss 0.00518254f
c50 40 Vss 7.20624e-19
c51 37 Vss 0.00663771f
c52 33 Vss 0.00663771f
c53 23 Vss 2.32346e-19
c54 20 Vss 0.211796f
c55 17 Vss 0.12596f
c56 15 Vss 0.0247918f
c57 4 Vss 0.137276f
r58 65 69 0.652036
r59 48 69 13.7956
r60 48 50 5.50157
r61 45 48 5.50157
r62 40 53 1.16709
r63 40 65 1.83386
r64 37 50 1.16709
r65 33 45 1.16709
r66 23 53 0.0476429
r67 21 23 0.326018
r68 21 23 0.1167
r69 20 24 0.652036
r70 20 23 6.7686
r71 17 53 0.357321
r72 15 23 0.326018
r73 15 17 0.40845
r74 8 37 0.185659
r75 6 33 0.185659
r76 4 24 3.8511
r77 2 17 3.44265
.ends

.subckt PM_G3_LATQ1_N2_GN 2 4 6 12 23 27 29 30 32 39 Vss
c44 39 Vss 0.0045172f
c45 32 Vss 8.57161e-19
c46 30 Vss 7.68504e-19
c47 29 Vss 0.00117249f
c48 27 Vss 0.00109299f
c49 23 Vss 0.00551775f
c50 12 Vss 0.171663f
c51 6 Vss 0.232172f
c52 4 Vss 0.00143442f
r53 32 39 1.16709
r54 29 32 0.531835
r55 29 30 1.70882
r56 25 30 0.652036
r57 25 27 4.91807
r58 23 27 1.16709
r59 14 39 0.197068
r60 12 16 0.652036
r61 12 14 4.668
r62 6 16 7.1187
r63 4 23 0.185659
r64 2 23 0.185659
.ends

.subckt PM_G3_LATQ1_N2_Q 2 4 13 18 Vss
c12 18 Vss 3.58669e-19
c13 13 Vss 0.004507f
c14 4 Vss 0.00143442f
r15 13 18 1.16709
r16 4 13 0.185659
r17 2 13 0.185659
.ends

.subckt PM_G3_LATQ1_N2_D 2 4 10 14 Vss
c14 14 Vss 4.15825e-19
c15 10 Vss 1.35847e-19
c16 2 Vss 0.475046f
r17 14 17 0.0416786
r18 10 17 1.16709
r19 4 10 7.7022
r20 2 10 7.7022
.ends

.subckt G3_LATQ1_N2  VDD VSS G Q D
*
* D	D
* Q	Q
* G	G
* VSS	VSS
* VDD	VDD
XI6.X0 N_GN_XI6.X0_D N_VSS_XI6.X0_PGD N_G_XI6.X0_CG N_VSS_XI6.X0_PGS
+ N_VDD_XI6.X0_S TIGFET_HPNW8
XI10.X0 N_Q_XI10.X0_D N_VDD_XI10.X0_PGD N_QN_XI10.X0_CG N_VDD_XI10.X0_PGS
+ N_VSS_XI10.X0_S TIGFET_HPNW8
XI9.X0 N_GN_XI9.X0_D N_VDD_XI9.X0_PGD N_G_XI9.X0_CG N_VDD_XI9.X0_PGS
+ N_VSS_XI9.X0_S TIGFET_HPNW8
XI8.X0 N_Q_XI8.X0_D N_VSS_XI8.X0_PGD N_QN_XI8.X0_CG N_VSS_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW8
XI11.X0 N_QN_XI11.X0_D N_VDD_XI11.X0_PGD N_D_XI11.X0_CG N_G_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW8
XI7.X0 N_QN_XI7.X0_D N_VSS_XI7.X0_PGD N_D_XI7.X0_CG N_GN_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW8
*
x_PM_G3_LATQ1_N2_VDD N_VDD_XI6.X0_S N_VDD_XI10.X0_PGD N_VDD_XI10.X0_PGS
+ N_VDD_XI9.X0_PGD N_VDD_XI9.X0_PGS N_VDD_XI8.X0_S N_VDD_XI11.X0_PGD
+ N_VDD_XI7.X0_S N_VDD_c_9_p N_VDD_c_5_p N_VDD_c_81_p N_VDD_c_15_p N_VDD_c_13_p
+ N_VDD_c_11_p N_VDD_c_7_p N_VDD_c_14_p N_VDD_c_6_p N_VDD_c_42_p N_VDD_c_19_p
+ N_VDD_c_46_p N_VDD_c_24_p N_VDD_c_10_p N_VDD_c_22_p N_VDD_c_12_p N_VDD_c_45_p
+ VDD N_VDD_c_27_p N_VDD_c_23_p Vss PM_G3_LATQ1_N2_VDD
x_PM_G3_LATQ1_N2_VSS N_VSS_XI6.X0_PGD N_VSS_XI6.X0_PGS N_VSS_XI10.X0_S
+ N_VSS_XI9.X0_S N_VSS_XI8.X0_PGD N_VSS_XI8.X0_PGS N_VSS_XI11.X0_S
+ N_VSS_XI7.X0_PGD N_VSS_c_94_n N_VSS_c_96_n N_VSS_c_139_p N_VSS_c_98_n
+ N_VSS_c_100_n N_VSS_c_102_n N_VSS_c_104_n N_VSS_c_106_n N_VSS_c_109_n
+ N_VSS_c_113_n N_VSS_c_117_n N_VSS_c_119_n N_VSS_c_123_n N_VSS_c_127_n
+ N_VSS_c_129_n N_VSS_c_130_n N_VSS_c_131_n N_VSS_c_132_n N_VSS_c_135_n
+ N_VSS_c_136_n N_VSS_c_137_n N_VSS_c_138_n VSS Vss PM_G3_LATQ1_N2_VSS
x_PM_G3_LATQ1_N2_G N_G_XI6.X0_CG N_G_XI9.X0_CG N_G_XI11.X0_PGS N_G_c_176_n
+ N_G_c_172_n N_G_c_173_n G N_G_c_175_n Vss PM_G3_LATQ1_N2_G
x_PM_G3_LATQ1_N2_QN N_QN_XI10.X0_CG N_QN_XI8.X0_CG N_QN_XI11.X0_D N_QN_XI7.X0_D
+ N_QN_c_197_n N_QN_c_198_n N_QN_c_214_n N_QN_c_199_n N_QN_c_201_n N_QN_c_204_n
+ N_QN_c_206_n N_QN_c_209_n N_QN_c_212_n Vss PM_G3_LATQ1_N2_QN
x_PM_G3_LATQ1_N2_GN N_GN_XI6.X0_D N_GN_XI9.X0_D N_GN_XI7.X0_PGS N_GN_c_243_n
+ N_GN_c_246_n N_GN_c_249_n N_GN_c_269_n N_GN_c_275_n N_GN_c_276_n N_GN_c_253_n
+ Vss PM_G3_LATQ1_N2_GN
x_PM_G3_LATQ1_N2_Q N_Q_XI10.X0_D N_Q_XI8.X0_D N_Q_c_287_n Q Vss PM_G3_LATQ1_N2_Q
x_PM_G3_LATQ1_N2_D N_D_XI11.X0_CG N_D_XI7.X0_CG N_D_c_304_n D Vss
+ PM_G3_LATQ1_N2_D
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI6.X0_PGD 0.00203852f
cc_2 N_VDD_XI10.X0_PGS N_VSS_XI6.X0_PGS 2.37403e-19
cc_3 N_VDD_XI10.X0_PGD N_VSS_XI8.X0_PGD 0.00203076f
cc_4 N_VDD_XI11.X0_PGD N_VSS_XI7.X0_PGD 2.37403e-19
cc_5 N_VDD_c_5_p N_VSS_c_94_n 0.00203852f
cc_6 N_VDD_c_6_p N_VSS_c_94_n 3.9313e-19
cc_7 N_VDD_c_7_p N_VSS_c_96_n 3.80615e-19
cc_8 N_VDD_c_6_p N_VSS_c_96_n 3.9313e-19
cc_9 N_VDD_c_9_p N_VSS_c_98_n 0.00203076f
cc_10 N_VDD_c_10_p N_VSS_c_98_n 2.95583e-19
cc_11 N_VDD_c_11_p N_VSS_c_100_n 2.64155e-19
cc_12 N_VDD_c_12_p N_VSS_c_100_n 8.58125e-19
cc_13 N_VDD_c_13_p N_VSS_c_102_n 2.12761e-19
cc_14 N_VDD_c_14_p N_VSS_c_102_n 9.5668e-19
cc_15 N_VDD_c_15_p N_VSS_c_104_n 2.64155e-19
cc_16 N_VDD_c_11_p N_VSS_c_104_n 2.69828e-19
cc_17 N_VDD_c_7_p N_VSS_c_106_n 4.61436e-19
cc_18 N_VDD_c_14_p N_VSS_c_106_n 0.00165395f
cc_19 N_VDD_c_19_p N_VSS_c_106_n 4.5625e-19
cc_20 N_VDD_c_7_p N_VSS_c_109_n 9.31121e-19
cc_21 N_VDD_c_6_p N_VSS_c_109_n 0.00161703f
cc_22 N_VDD_c_22_p N_VSS_c_109_n 7.09654e-19
cc_23 N_VDD_c_23_p N_VSS_c_109_n 3.48267e-19
cc_24 N_VDD_c_24_p N_VSS_c_113_n 9.52068e-19
cc_25 N_VDD_c_10_p N_VSS_c_113_n 0.00141228f
cc_26 N_VDD_c_12_p N_VSS_c_113_n 0.00257912f
cc_27 N_VDD_c_27_p N_VSS_c_113_n 3.48267e-19
cc_28 N_VDD_c_7_p N_VSS_c_117_n 2.12713e-19
cc_29 N_VDD_c_22_p N_VSS_c_117_n 8.43845e-19
cc_30 N_VDD_c_7_p N_VSS_c_119_n 4.24454e-19
cc_31 N_VDD_c_6_p N_VSS_c_119_n 2.26455e-19
cc_32 N_VDD_c_22_p N_VSS_c_119_n 3.84769e-19
cc_33 N_VDD_c_23_p N_VSS_c_119_n 6.489e-19
cc_34 N_VDD_c_24_p N_VSS_c_123_n 3.82294e-19
cc_35 N_VDD_c_10_p N_VSS_c_123_n 0.00114511f
cc_36 N_VDD_c_12_p N_VSS_c_123_n 9.55109e-19
cc_37 N_VDD_c_27_p N_VSS_c_123_n 6.46219e-19
cc_38 N_VDD_c_7_p N_VSS_c_127_n 0.00468852f
cc_39 N_VDD_c_14_p N_VSS_c_127_n 0.00657271f
cc_40 N_VDD_c_14_p N_VSS_c_129_n 0.00377187f
cc_41 N_VDD_c_6_p N_VSS_c_130_n 0.00345737f
cc_42 N_VDD_c_42_p N_VSS_c_131_n 0.00106538f
cc_43 N_VDD_c_19_p N_VSS_c_132_n 0.00353938f
cc_44 N_VDD_c_10_p N_VSS_c_132_n 0.00581493f
cc_45 N_VDD_c_45_p N_VSS_c_132_n 9.99051e-19
cc_46 N_VDD_c_46_p N_VSS_c_135_n 0.0010616f
cc_47 N_VDD_c_6_p N_VSS_c_136_n 0.00566938f
cc_48 N_VDD_c_14_p N_VSS_c_137_n 9.16632e-19
cc_49 N_VDD_c_6_p N_VSS_c_138_n 7.74609e-19
cc_50 N_VDD_c_15_p N_G_XI11.X0_PGS 0.00163289f
cc_51 N_VDD_XI9.X0_PGD N_G_c_172_n 3.96934e-19
cc_52 N_VDD_XI9.X0_PGS N_G_c_173_n 4.08222e-19
cc_53 N_VDD_c_14_p G 5.04211e-19
cc_54 N_VDD_c_14_p N_G_c_175_n 5.56409e-19
cc_55 N_VDD_XI10.X0_PGD N_QN_c_197_n 4.07423e-19
cc_56 N_VDD_c_27_p N_QN_c_198_n 0.00100159f
cc_57 N_VDD_c_11_p N_QN_c_199_n 3.43419e-19
cc_58 N_VDD_c_12_p N_QN_c_199_n 3.48267e-19
cc_59 N_VDD_c_14_p N_QN_c_201_n 4.08289e-19
cc_60 N_VDD_c_24_p N_QN_c_201_n 2.98644e-19
cc_61 N_VDD_c_27_p N_QN_c_201_n 3.15998e-19
cc_62 N_VDD_c_11_p N_QN_c_204_n 3.48267e-19
cc_63 N_VDD_c_12_p N_QN_c_204_n 9.04108e-19
cc_64 N_VDD_c_6_p N_QN_c_206_n 3.90695e-19
cc_65 N_VDD_c_10_p N_QN_c_206_n 3.49463e-19
cc_66 N_VDD_c_12_p N_QN_c_206_n 3.67848e-19
cc_67 N_VDD_c_14_p N_QN_c_209_n 6.60137e-19
cc_68 N_VDD_c_24_p N_QN_c_209_n 3.43988e-19
cc_69 N_VDD_c_27_p N_QN_c_209_n 2.68747e-19
cc_70 N_VDD_c_14_p N_QN_c_212_n 3.90734e-19
cc_71 N_VDD_XI9.X0_PGS N_GN_c_243_n 3.40745e-19
cc_72 N_VDD_c_15_p N_GN_c_243_n 2.49684e-19
cc_73 N_VDD_c_11_p N_GN_c_243_n 3.08361e-19
cc_74 N_VDD_c_13_p N_GN_c_246_n 3.43419e-19
cc_75 N_VDD_c_7_p N_GN_c_246_n 3.72199e-19
cc_76 N_VDD_c_6_p N_GN_c_246_n 3.4118e-19
cc_77 N_VDD_c_13_p N_GN_c_249_n 3.48267e-19
cc_78 N_VDD_c_7_p N_GN_c_249_n 7.94301e-19
cc_79 N_VDD_c_14_p N_GN_c_249_n 0.0010243f
cc_80 N_VDD_c_6_p N_GN_c_249_n 4.77682e-19
cc_81 N_VDD_c_81_p N_GN_c_253_n 3.88849e-19
cc_82 N_VDD_c_22_p N_GN_c_253_n 2.02851e-19
cc_83 N_VDD_c_11_p N_Q_c_287_n 3.43419e-19
cc_84 N_VDD_c_10_p N_Q_c_287_n 3.4118e-19
cc_85 N_VDD_c_12_p N_Q_c_287_n 3.48267e-19
cc_86 N_VDD_c_11_p Q 3.48267e-19
cc_87 N_VDD_c_10_p Q 4.58391e-19
cc_88 N_VDD_c_12_p Q 7.09569e-19
cc_89 N_VDD_c_15_p N_D_XI11.X0_CG 4.20341e-19
cc_90 N_VSS_c_139_p N_G_c_176_n 9.37683e-19
cc_91 N_VSS_XI6.X0_PGD N_G_c_172_n 4.04227e-19
cc_92 N_VSS_c_109_n G 3.00355e-19
cc_93 N_VSS_c_119_n G 3.2351e-19
cc_94 N_VSS_c_127_n G 2.86445e-19
cc_95 N_VSS_c_109_n N_G_c_175_n 3.2351e-19
cc_96 N_VSS_c_119_n N_G_c_175_n 2.68747e-19
cc_97 N_VSS_XI8.X0_PGD N_QN_c_197_n 3.93738e-19
cc_98 N_VSS_c_104_n N_QN_c_214_n 3.43419e-19
cc_99 N_VSS_c_117_n N_QN_c_214_n 3.48267e-19
cc_100 N_VSS_c_132_n N_QN_c_201_n 2.32769e-19
cc_101 N_VSS_c_104_n N_QN_c_204_n 3.48267e-19
cc_102 N_VSS_c_117_n N_QN_c_204_n 8.62542e-19
cc_103 N_VSS_c_113_n N_QN_c_206_n 2.72578e-19
cc_104 N_VSS_c_117_n N_QN_c_206_n 6.59201e-19
cc_105 N_VSS_c_132_n N_QN_c_206_n 5.73383e-19
cc_106 N_VSS_c_136_n N_QN_c_206_n 7.86339e-19
cc_107 N_VSS_c_109_n N_QN_c_212_n 4.50267e-19
cc_108 N_VSS_c_127_n N_QN_c_212_n 0.00182171f
cc_109 N_VSS_c_100_n N_GN_XI7.X0_PGS 0.00172633f
cc_110 N_VSS_XI8.X0_PGS N_GN_c_243_n 6.82193e-19
cc_111 N_VSS_c_104_n N_GN_c_246_n 3.43419e-19
cc_112 N_VSS_c_117_n N_GN_c_246_n 3.48267e-19
cc_113 N_VSS_c_104_n N_GN_c_249_n 3.48267e-19
cc_114 N_VSS_c_117_n N_GN_c_249_n 4.99861e-19
cc_115 N_VSS_c_127_n N_GN_c_249_n 5.59824e-19
cc_116 N_VSS_c_113_n N_GN_c_253_n 2.02167e-19
cc_117 N_VSS_c_123_n N_GN_c_253_n 3.56129e-19
cc_118 N_VSS_c_102_n N_Q_c_287_n 3.43419e-19
cc_119 N_VSS_c_106_n N_Q_c_287_n 3.48267e-19
cc_120 N_VSS_c_106_n Q 8.15956e-19
cc_121 N_VSS_c_100_n N_D_XI11.X0_CG 4.20341e-19
cc_122 N_G_c_172_n N_QN_c_197_n 0.00398811f
cc_123 G N_QN_c_201_n 4.48861e-19
cc_124 N_G_c_175_n N_QN_c_201_n 4.54925e-19
cc_125 G N_QN_c_209_n 4.56568e-19
cc_126 N_G_c_175_n N_QN_c_209_n 0.00268575f
cc_127 N_G_c_173_n N_GN_c_243_n 0.00842907f
cc_128 N_G_c_172_n N_GN_c_246_n 6.8653e-19
cc_129 N_G_c_172_n N_GN_c_249_n 3.82175e-19
cc_130 G N_GN_c_249_n 0.00151253f
cc_131 N_G_c_175_n N_GN_c_249_n 9.72448e-19
cc_132 N_G_c_172_n N_GN_c_269_n 3.75306e-19
cc_133 N_G_c_172_n N_GN_c_253_n 0.00395135f
cc_134 N_G_c_175_n N_GN_c_253_n 2.41671e-19
cc_135 N_G_XI11.X0_PGS N_D_XI11.X0_CG 0.00435077f
cc_136 N_QN_c_197_n N_GN_XI7.X0_PGS 0.00196434f
cc_137 N_QN_c_204_n N_GN_c_249_n 0.0010213f
cc_138 N_QN_c_206_n N_GN_c_269_n 9.45997e-19
cc_139 N_QN_c_206_n N_GN_c_275_n 0.00125885f
cc_140 N_QN_c_206_n N_GN_c_276_n 9.71021e-19
cc_141 N_QN_c_197_n N_GN_c_253_n 0.00340055f
cc_142 N_QN_c_209_n N_GN_c_253_n 2.75519e-19
cc_143 N_QN_c_197_n N_Q_c_287_n 6.8653e-19
cc_144 N_QN_c_197_n N_D_XI11.X0_CG 3.26559e-19
cc_145 N_QN_c_204_n N_D_XI11.X0_CG 0.0010503f
cc_146 N_QN_c_204_n N_D_c_304_n 0.00130556f
cc_147 N_QN_c_204_n D 0.00141415f
cc_148 N_QN_c_206_n D 0.00146947f
cc_149 N_GN_c_275_n N_Q_c_287_n 4.09054e-19
cc_150 N_GN_c_275_n Q 5.11868e-19
cc_151 N_GN_XI7.X0_PGS N_D_XI11.X0_CG 0.0048787f
cc_152 N_GN_c_243_n N_D_c_304_n 0.00333193f
cc_153 N_GN_c_276_n N_D_c_304_n 3.73302e-19
cc_154 N_GN_c_253_n N_D_c_304_n 8.5422e-19
cc_155 N_GN_c_276_n D 2.85187e-19
cc_156 N_GN_c_253_n D 3.48267e-19
*
.ends
*
*
.subckt LATQ1_HPNW8 D G Q VDD VSS
xgate (VDD VSS G Q D) G3_LATQ1_N2
.ends
*
* File: G4_MAJ3_N2.pex.netlist
* Created: Fri Mar  4 11:26:54 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MAJ3_N2_VDD 2 4 7 11 27 28 30 31 32 44 48 52 54 56 57 58 61 63 67
+ 69 70 73 77 79 80 90 95 Vss
c77 95 Vss 0.00486523f
c78 90 Vss 0.00461066f
c79 80 Vss 4.52364e-19
c80 79 Vss 4.28405e-19
c81 77 Vss 4.66438e-19
c82 73 Vss 8.57616e-19
c83 70 Vss 8.64091e-19
c84 69 Vss 0.00558016f
c85 67 Vss 0.00139758f
c86 63 Vss 0.00140124f
c87 58 Vss 8.64091e-19
c88 57 Vss 0.00559492f
c89 56 Vss 0.00209681f
c90 54 Vss 0.00571364f
c91 52 Vss 0.00207954f
c92 48 Vss 0.00382489f
c93 44 Vss 0.00532438f
c94 32 Vss 0.035607f
c95 31 Vss 0.100823f
c96 28 Vss 0.035607f
c97 27 Vss 0.100961f
c98 11 Vss 0.266772f
c99 7 Vss 0.268336f
r100 77 95 1.16709
r101 75 77 2.16729
r102 73 90 1.16709
r103 71 73 2.16729
r104 69 75 0.652036
r105 69 70 10.1279
r106 65 80 0.0828784
r107 65 67 1.82344
r108 61 63 1.167
r109 59 79 0.0828784
r110 59 61 0.656438
r111 57 71 0.652036
r112 57 58 10.1279
r113 56 70 0.652036
r114 55 80 0.551426
r115 55 56 4.58464
r116 54 80 0.551426
r117 53 79 0.551426
r118 53 54 9.66943
r119 52 79 0.551426
r120 51 58 0.652036
r121 51 52 4.58464
r122 48 67 1.16709
r123 44 63 1.16709
r124 34 95 0.0476429
r125 32 34 1.45875
r126 31 38 0.652036
r127 31 34 1.45875
r128 30 90 0.0476429
r129 28 30 1.45875
r130 27 35 0.652036
r131 27 30 1.45875
r132 24 32 0.652036
r133 21 28 0.652036
r134 11 38 3.8511
r135 11 24 3.8511
r136 7 35 3.8511
r137 7 21 3.8511
r138 4 48 0.185659
r139 2 44 0.185659
.ends

.subckt PM_G4_MAJ3_N2_VSS 3 7 10 12 27 28 30 31 32 45 49 52 57 62 67 70 73 78 91
+ 92 93 94 95 104 114 115 117 Vss
c83 115 Vss 3.75522e-19
c84 114 Vss 3.75522e-19
c85 110 Vss 0.00128107f
c86 104 Vss 0.00335813f
c87 95 Vss 8.27105e-19
c88 94 Vss 0.00156442f
c89 93 Vss 8.27105e-19
c90 92 Vss 0.00156442f
c91 91 Vss 0.00686995f
c92 78 Vss 0.00393332f
c93 73 Vss 0.00431768f
c94 70 Vss 0.00351391f
c95 67 Vss 0.00277973f
c96 62 Vss 0.00186148f
c97 57 Vss 0.00131291f
c98 52 Vss 0.00112626f
c99 49 Vss 0.00527641f
c100 45 Vss 0.00377692f
c101 32 Vss 0.0350852f
c102 31 Vss 0.0994129f
c103 30 Vss 9.50876e-20
c104 28 Vss 0.0350852f
c105 27 Vss 0.0994129f
c106 7 Vss 0.267138f
c107 3 Vss 0.268863f
r108 110 117 0.326018
r109 106 115 0.494161
r110 105 114 0.494161
r111 104 117 0.326018
r112 104 105 7.46046
r113 100 115 0.128424
r114 96 114 0.128424
r115 94 115 0.494161
r116 94 95 4.37625
r117 92 114 0.494161
r118 92 93 4.37625
r119 91 95 0.652036
r120 90 93 0.652036
r121 90 91 21.5061
r122 70 106 8.04396
r123 67 70 5.835
r124 62 110 5.2515
r125 57 78 1.16709
r126 57 100 2.16729
r127 52 73 1.16709
r128 52 96 2.16729
r129 49 67 1.16709
r130 45 62 1.16709
r131 34 78 0.0476429
r132 32 34 1.45875
r133 31 38 0.652036
r134 31 34 1.45875
r135 30 73 0.0476429
r136 28 30 1.45875
r137 27 35 0.652036
r138 27 30 1.45875
r139 24 32 0.652036
r140 21 28 0.652036
r141 12 49 0.185659
r142 10 45 0.185659
r143 7 38 3.8511
r144 7 24 3.8511
r145 3 35 3.8511
r146 3 21 3.8511
.ends

.subckt PM_G4_MAJ3_N2_A 1 2 4 6 9 13 31 53 57 62 67 71 74 76 78 81 89 91 99 100
+ 102 111 Vss
c78 111 Vss 0.00528881f
c79 102 Vss 0.00500597f
c80 99 Vss 0.00422425f
c81 96 Vss 7.53731e-19
c82 91 Vss 7.84512e-19
c83 89 Vss 8.92851e-19
c84 85 Vss 0.00253152f
c85 81 Vss 7.20282e-19
c86 78 Vss 0.0011176f
c87 77 Vss 0.00146569f
c88 76 Vss 0.00441934f
c89 71 Vss 0.00722904f
c90 67 Vss 0.00399277f
c91 62 Vss 0.00496845f
c92 57 Vss 0.135055f
c93 53 Vss 0.12803f
c94 31 Vss 0.215113f
c95 27 Vss 0.126125f
c96 25 Vss 0.0247918f
c97 9 Vss 1.22732f
c98 2 Vss 0.139046f
r99 111 114 0.1
r100 98 111 1.16709
r101 98 100 0.490235
r102 98 99 0.490235
r103 94 102 1.16709
r104 91 94 1.08364
r105 87 89 2.50071
r106 85 87 0.653045
r107 85 100 1.5949
r108 84 96 0.466409
r109 84 99 6.9631
r110 79 96 0.152298
r111 79 81 2.50071
r112 77 96 0.466409
r113 77 78 1.7116
r114 75 78 0.653045
r115 75 76 8.7525
r116 72 91 0.0685365
r117 72 74 1.45875
r118 71 76 0.652036
r119 71 74 8.7525
r120 67 89 1.16709
r121 62 81 1.16709
r122 55 57 4.53833
r123 52 114 0.0238214
r124 52 53 2.26917
r125 49 52 2.26917
r126 44 57 0.00605528
r127 43 53 0.00605528
r128 40 55 0.00605528
r129 39 49 0.00605528
r130 34 102 0.0476429
r131 32 34 0.326018
r132 32 34 0.1167
r133 31 35 0.652036
r134 31 34 6.7686
r135 27 102 0.357321
r136 25 34 0.326018
r137 25 27 0.40845
r138 13 44 3.8511
r139 13 40 3.8511
r140 9 13 15.4044
r141 9 43 3.8511
r142 9 13 15.4044
r143 9 39 3.8511
r144 6 67 0.185659
r145 4 62 0.185659
r146 2 35 3.8511
r147 1 27 3.44265
.ends

.subckt PM_G4_MAJ3_N2_BI 2 4 5 6 20 29 34 39 44 54 59 68 74 75 83 Vss
c58 83 Vss 4.27892e-19
c59 75 Vss 3.15444e-19
c60 74 Vss 7.27663e-19
c61 68 Vss 0.00155105f
c62 59 Vss 0.00147096f
c63 54 Vss 0.00139826f
c64 44 Vss 0.00152385f
c65 39 Vss 0.00577944f
c66 34 Vss 0.00175738f
c67 29 Vss 0.00439389f
c68 20 Vss 0.111942f
c69 5 Vss 0.111942f
c70 4 Vss 0.00143442f
r71 79 83 0.655813
r72 74 75 0.65228
r73 73 74 3.42052
r74 68 73 0.65409
r75 44 59 1.16709
r76 44 75 2.1395
r77 39 54 1.16709
r78 39 83 12.0712
r79 39 68 1.96931
r80 34 51 1.16709
r81 34 79 2.334
r82 29 51 0.1
r83 20 59 0.50025
r84 17 54 0.50025
r85 6 20 3.09255
r86 5 17 3.09255
r87 4 29 0.185659
r88 2 29 0.185659
.ends

.subckt PM_G4_MAJ3_N2_AI 2 4 7 11 31 37 43 46 51 60 69 Vss
c44 69 Vss 4.10597e-19
c45 60 Vss 0.00527726f
c46 51 Vss 0.00584502f
c47 46 Vss 0.00110084f
c48 43 Vss 0.00447686f
c49 37 Vss 0.127877f
c50 31 Vss 0.134503f
c51 7 Vss 1.21876f
c52 4 Vss 0.00143442f
r53 65 69 0.652036
r54 60 63 0.1
r55 51 63 1.16709
r56 51 69 13.7539
r57 46 65 2.58407
r58 43 46 1.16709
r59 36 60 0.0238214
r60 36 37 2.334
r61 33 36 2.20433
r62 29 31 4.53833
r63 26 37 0.00605528
r64 25 31 0.00605528
r65 22 33 0.00605528
r66 21 29 0.00605528
r67 11 26 3.8511
r68 11 22 3.8511
r69 7 11 15.4044
r70 7 25 3.8511
r71 7 11 15.4044
r72 7 21 3.8511
r73 4 43 0.185659
r74 2 43 0.185659
.ends

.subckt PM_G4_MAJ3_N2_B 1 2 3 4 13 14 24 42 46 49 54 59 64 69 77 78 84 91 96 97
+ Vss
c68 97 Vss 4.67818e-19
c69 96 Vss 0.00212566f
c70 91 Vss 9.32419e-19
c71 84 Vss 5.17496e-19
c72 78 Vss 3.17701e-19
c73 77 Vss 0.00357974f
c74 69 Vss 0.00148026f
c75 64 Vss 0.0010348f
c76 59 Vss 0.00464385f
c77 54 Vss 0.00163559f
c78 49 Vss 7.01001e-19
c79 46 Vss 5.25457e-19
c80 42 Vss 5.46753e-19
c81 24 Vss 0.111942f
c82 17 Vss 0.0247918f
c83 14 Vss 0.0349292f
c84 13 Vss 0.183407f
c85 4 Vss 0.111942f
c86 2 Vss 0.111095f
c87 1 Vss 0.118069f
r88 95 97 0.65409
r89 95 96 3.42052
r90 91 96 0.65228
r91 87 91 2.1006
r92 84 87 2.04225
r93 77 84 0.0685365
r94 77 78 10.3363
r95 73 78 0.652036
r96 54 69 1.16709
r97 54 97 2.00578
r98 49 64 1.16709
r99 49 87 0.0416786
r100 42 59 1.16709
r101 42 73 2.16729
r102 42 46 0.0530455
r103 36 59 0.238214
r104 33 69 0.50025
r105 24 64 0.50025
r106 22 36 0.262036
r107 17 36 0.326018
r108 17 22 0.05835
r109 14 36 6.7686
r110 13 36 0.326018
r111 13 36 0.1167
r112 9 14 0.652036
r113 4 33 3.09255
r114 3 24 3.09255
r115 2 22 3.09255
r116 1 9 3.1509
.ends

.subckt PM_G4_MAJ3_N2_C 2 4 12 17 20 25 51 Vss
c18 25 Vss 0.00550018f
c19 20 Vss 7.32915e-19
c20 17 Vss 0.00502472f
c21 12 Vss 0.00387713f
r22 25 51 1.78697
r23 20 51 8.27841
r24 17 25 1.16709
r25 12 20 1.16709
r26 4 17 0.185659
r27 2 12 0.185659
.ends

.subckt PM_G4_MAJ3_N2_Z 2 4 6 8 23 27 30 33 Vss
c30 30 Vss 0.00298505f
c31 27 Vss 0.00857889f
c32 23 Vss 0.00745393f
c33 8 Vss 0.00143442f
c34 6 Vss 0.00143442f
r35 33 35 6.04339
r36 30 33 4.95975
r37 27 35 1.16709
r38 23 30 1.16709
r39 8 27 0.185659
r40 6 23 0.185659
r41 4 27 0.185659
r42 2 23 0.185659
.ends

.subckt G4_MAJ3_N2  VDD VSS A B C Z
*
* Z	Z
* C	C
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI11.X0 N_BI_XI11.X0_D N_VSS_XI11.X0_PGD N_B_XI11.X0_CG N_VSS_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW8
XI10.X0 N_AI_XI10.X0_D N_VSS_XI10.X0_PGD N_A_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW8
XI9.X0 N_BI_XI9.X0_D N_VDD_XI9.X0_PGD N_B_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW8
XI0.X0 N_AI_XI0.X0_D N_VDD_XI0.X0_PGD N_A_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_AI_XI15.X0_PGD N_BI_XI15.X0_CG N_AI_XI15.X0_PGD
+ N_A_XI15.X0_S TIGFET_HPNW8
XI13.X0 N_Z_XI13.X0_D N_AI_XI13.X0_PGD N_B_XI13.X0_CG N_AI_XI13.X0_PGD
+ N_C_XI13.X0_S TIGFET_HPNW8
XI14.X0 N_Z_XI14.X0_D N_A_XI14.X0_PGD N_B_XI14.X0_CG N_A_XI14.X0_PGD
+ N_A_XI14.X0_S TIGFET_HPNW8
XI12.X0 N_Z_XI12.X0_D N_A_XI12.X0_PGD N_BI_XI12.X0_CG N_A_XI12.X0_PGD
+ N_C_XI12.X0_S TIGFET_HPNW8
*
x_PM_G4_MAJ3_N2_VDD N_VDD_XI11.X0_S N_VDD_XI10.X0_S N_VDD_XI9.X0_PGD
+ N_VDD_XI0.X0_PGD N_VDD_c_62_p N_VDD_c_4_p N_VDD_c_72_p N_VDD_c_63_p
+ N_VDD_c_8_p N_VDD_c_55_p N_VDD_c_64_p N_VDD_c_6_p N_VDD_c_32_p N_VDD_c_3_p
+ N_VDD_c_5_p N_VDD_c_38_p VDD N_VDD_c_37_p N_VDD_c_39_p N_VDD_c_9_p
+ N_VDD_c_41_p N_VDD_c_13_p N_VDD_c_17_p N_VDD_c_34_p N_VDD_c_35_p N_VDD_c_14_p
+ N_VDD_c_18_p Vss PM_G4_MAJ3_N2_VDD
x_PM_G4_MAJ3_N2_VSS N_VSS_XI11.X0_PGD N_VSS_XI10.X0_PGD N_VSS_XI9.X0_S
+ N_VSS_XI0.X0_S N_VSS_c_81_n N_VSS_c_83_n N_VSS_c_135_p N_VSS_c_85_n
+ N_VSS_c_87_n N_VSS_c_123_p N_VSS_c_125_p N_VSS_c_88_n N_VSS_c_92_n
+ N_VSS_c_96_n N_VSS_c_97_n N_VSS_c_100_n N_VSS_c_101_n N_VSS_c_105_n
+ N_VSS_c_108_n N_VSS_c_113_n N_VSS_c_115_n N_VSS_c_116_n N_VSS_c_118_n
+ N_VSS_c_119_n N_VSS_c_120_n N_VSS_c_121_n VSS Vss PM_G4_MAJ3_N2_VSS
x_PM_G4_MAJ3_N2_A N_A_XI10.X0_CG N_A_XI0.X0_CG N_A_XI15.X0_S N_A_XI14.X0_S
+ N_A_XI14.X0_PGD N_A_XI12.X0_PGD N_A_c_161_n N_A_c_201_p N_A_c_203_p
+ N_A_c_172_n N_A_c_228_p N_A_c_162_n A N_A_c_179_n N_A_c_167_n N_A_c_223_p
+ N_A_c_230_p N_A_c_169_n N_A_c_187_p N_A_c_215_p N_A_c_170_n N_A_c_216_p Vss
+ PM_G4_MAJ3_N2_A
x_PM_G4_MAJ3_N2_BI N_BI_XI11.X0_D N_BI_XI9.X0_D N_BI_XI15.X0_CG N_BI_XI12.X0_CG
+ N_BI_c_252_n N_BI_c_239_n N_BI_c_241_n N_BI_c_249_n N_BI_c_257_n N_BI_c_258_n
+ N_BI_c_259_n N_BI_c_260_n N_BI_c_280_p N_BI_c_283_p N_BI_c_261_n Vss
+ PM_G4_MAJ3_N2_BI
x_PM_G4_MAJ3_N2_AI N_AI_XI10.X0_D N_AI_XI0.X0_D N_AI_XI15.X0_PGD
+ N_AI_XI13.X0_PGD N_AI_c_299_n N_AI_c_300_n N_AI_c_301_n N_AI_c_303_n
+ N_AI_c_306_n N_AI_c_315_n N_AI_c_316_n Vss PM_G4_MAJ3_N2_AI
x_PM_G4_MAJ3_N2_B N_B_XI11.X0_CG N_B_XI9.X0_CG N_B_XI13.X0_CG N_B_XI14.X0_CG
+ N_B_c_341_n N_B_c_355_n N_B_c_393_n N_B_c_342_n B N_B_c_374_n N_B_c_359_n
+ N_B_c_346_n N_B_c_378_n N_B_c_364_n N_B_c_351_n N_B_c_370_n N_B_c_371_n
+ N_B_c_387_n N_B_c_390_n N_B_c_391_n Vss PM_G4_MAJ3_N2_B
x_PM_G4_MAJ3_N2_C N_C_XI13.X0_S N_C_XI12.X0_S N_C_c_409_n N_C_c_422_p
+ N_C_c_410_n N_C_c_412_n C Vss PM_G4_MAJ3_N2_C
x_PM_G4_MAJ3_N2_Z N_Z_XI15.X0_D N_Z_XI13.X0_D N_Z_XI14.X0_D N_Z_XI12.X0_D
+ N_Z_c_427_n N_Z_c_451_n N_Z_c_432_n Z Vss PM_G4_MAJ3_N2_Z
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI11.X0_PGD 0.00200884f
cc_2 N_VDD_XI0.X0_PGD N_VSS_XI10.X0_PGD 0.0020057f
cc_3 N_VDD_c_3_p N_VSS_XI10.X0_PGD 2.76462e-19
cc_4 N_VDD_c_4_p N_VSS_c_81_n 0.00200884f
cc_5 N_VDD_c_5_p N_VSS_c_81_n 3.23379e-19
cc_6 N_VDD_c_6_p N_VSS_c_83_n 2.76462e-19
cc_7 N_VDD_c_5_p N_VSS_c_83_n 3.9313e-19
cc_8 N_VDD_c_8_p N_VSS_c_85_n 0.0020057f
cc_9 N_VDD_c_9_p N_VSS_c_85_n 2.84318e-19
cc_10 N_VDD_c_9_p N_VSS_c_87_n 3.9313e-19
cc_11 N_VDD_c_6_p N_VSS_c_88_n 4.35319e-19
cc_12 N_VDD_c_5_p N_VSS_c_88_n 0.00161703f
cc_13 N_VDD_c_13_p N_VSS_c_88_n 9.22325e-19
cc_14 N_VDD_c_14_p N_VSS_c_88_n 3.48267e-19
cc_15 N_VDD_c_3_p N_VSS_c_92_n 4.76491e-19
cc_16 N_VDD_c_9_p N_VSS_c_92_n 0.00161703f
cc_17 N_VDD_c_17_p N_VSS_c_92_n 8.59637e-19
cc_18 N_VDD_c_18_p N_VSS_c_92_n 3.48267e-19
cc_19 N_VDD_c_13_p N_VSS_c_96_n 8.49247e-19
cc_20 N_VDD_XI0.X0_PGD N_VSS_c_97_n 2.8629e-19
cc_21 N_VDD_c_17_p N_VSS_c_97_n 0.00515616f
cc_22 N_VDD_c_18_p N_VSS_c_97_n 9.58524e-19
cc_23 N_VDD_c_9_p N_VSS_c_100_n 0.00401341f
cc_24 N_VDD_c_6_p N_VSS_c_101_n 3.66936e-19
cc_25 N_VDD_c_5_p N_VSS_c_101_n 2.26455e-19
cc_26 N_VDD_c_13_p N_VSS_c_101_n 3.99794e-19
cc_27 N_VDD_c_14_p N_VSS_c_101_n 6.489e-19
cc_28 N_VDD_c_9_p N_VSS_c_105_n 2.26455e-19
cc_29 N_VDD_c_17_p N_VSS_c_105_n 3.99794e-19
cc_30 N_VDD_c_18_p N_VSS_c_105_n 6.489e-19
cc_31 N_VDD_c_6_p N_VSS_c_108_n 0.00335989f
cc_32 N_VDD_c_32_p N_VSS_c_108_n 0.00777551f
cc_33 N_VDD_c_3_p N_VSS_c_108_n 0.0031218f
cc_34 N_VDD_c_34_p N_VSS_c_108_n 0.00104624f
cc_35 N_VDD_c_35_p N_VSS_c_108_n 0.0010706f
cc_36 N_VDD_c_5_p N_VSS_c_113_n 0.00329944f
cc_37 N_VDD_c_37_p N_VSS_c_113_n 3.33664e-19
cc_38 N_VDD_c_38_p N_VSS_c_115_n 0.00106538f
cc_39 N_VDD_c_39_p N_VSS_c_116_n 3.33664e-19
cc_40 N_VDD_c_9_p N_VSS_c_116_n 0.00329944f
cc_41 N_VDD_c_41_p N_VSS_c_118_n 0.00106538f
cc_42 N_VDD_c_5_p N_VSS_c_119_n 0.00554732f
cc_43 N_VDD_c_5_p N_VSS_c_120_n 7.74609e-19
cc_44 N_VDD_c_9_p N_VSS_c_121_n 7.74609e-19
cc_45 N_VDD_XI0.X0_PGD N_A_c_161_n 3.94724e-19
cc_46 N_VDD_XI0.X0_PGD N_A_c_162_n 4.99274e-19
cc_47 N_VDD_c_5_p N_A_c_162_n 2.55296e-19
cc_48 N_VDD_c_9_p N_A_c_162_n 2.95925e-19
cc_49 N_VDD_c_17_p N_A_c_162_n 3.33497e-19
cc_50 N_VDD_c_18_p N_A_c_162_n 2.46105e-19
cc_51 N_VDD_c_13_p N_A_c_167_n 5.45771e-19
cc_52 N_VDD_c_14_p N_A_c_167_n 4.10732e-19
cc_53 N_VDD_c_32_p N_A_c_169_n 9.17955e-19
cc_54 N_VDD_c_32_p N_A_c_170_n 4.71221e-19
cc_55 N_VDD_c_55_p N_BI_c_239_n 3.43419e-19
cc_56 N_VDD_c_37_p N_BI_c_239_n 3.72199e-19
cc_57 N_VDD_c_55_p N_BI_c_241_n 3.48267e-19
cc_58 N_VDD_c_5_p N_BI_c_241_n 4.22613e-19
cc_59 N_VDD_c_37_p N_BI_c_241_n 5.2846e-19
cc_60 N_VDD_XI9.X0_PGD N_AI_XI15.X0_PGD 2.83823e-19
cc_61 N_VDD_XI0.X0_PGD N_AI_XI15.X0_PGD 3.10667e-19
cc_62 N_VDD_c_62_p N_AI_c_299_n 2.83823e-19
cc_63 N_VDD_c_63_p N_AI_c_300_n 3.10667e-19
cc_64 N_VDD_c_64_p N_AI_c_301_n 3.43419e-19
cc_65 N_VDD_c_39_p N_AI_c_301_n 3.72199e-19
cc_66 N_VDD_c_64_p N_AI_c_303_n 3.48267e-19
cc_67 N_VDD_c_39_p N_AI_c_303_n 5.226e-19
cc_68 N_VDD_c_9_p N_AI_c_303_n 4.34701e-19
cc_69 N_VDD_c_17_p N_AI_c_306_n 9.61607e-19
cc_70 N_VDD_XI9.X0_PGD N_B_c_341_n 3.99218e-19
cc_71 N_VDD_c_32_p N_B_c_342_n 3.87456e-19
cc_72 N_VDD_c_72_p B 3.02565e-19
cc_73 N_VDD_c_13_p B 4.44319e-19
cc_74 N_VDD_c_14_p B 3.49905e-19
cc_75 N_VDD_c_13_p N_B_c_346_n 3.43988e-19
cc_76 N_VDD_c_14_p N_B_c_346_n 2.68747e-19
cc_77 N_VDD_c_18_p N_B_c_346_n 4.88234e-19
cc_78 N_VSS_XI10.X0_PGD N_A_c_161_n 3.91527e-19
cc_79 N_VSS_c_123_p N_A_c_172_n 3.43419e-19
cc_80 N_VSS_c_123_p N_A_c_162_n 2.69869e-19
cc_81 N_VSS_c_125_p N_A_c_162_n 5.38503e-19
cc_82 N_VSS_c_96_n N_A_c_162_n 3.16844e-19
cc_83 N_VSS_c_97_n N_A_c_162_n 8.92829e-19
cc_84 N_VSS_c_100_n N_A_c_162_n 2.86582e-19
cc_85 N_VSS_c_119_n N_A_c_162_n 2.99293e-19
cc_86 N_VSS_c_96_n N_A_c_179_n 0.00223349f
cc_87 N_VSS_c_96_n N_A_c_167_n 0.00150218f
cc_88 N_VSS_c_92_n N_A_c_169_n 3.34005e-19
cc_89 N_VSS_c_105_n N_A_c_169_n 6.63553e-19
cc_90 N_VSS_c_108_n N_A_c_169_n 5.04162e-19
cc_91 N_VSS_c_135_p N_A_c_170_n 2.02217e-19
cc_92 N_VSS_c_92_n N_A_c_170_n 3.2351e-19
cc_93 N_VSS_c_105_n N_A_c_170_n 2.68747e-19
cc_94 N_VSS_c_123_p N_BI_c_239_n 3.43419e-19
cc_95 N_VSS_c_123_p N_BI_c_241_n 3.48267e-19
cc_96 N_VSS_c_96_n N_BI_c_241_n 0.00105024f
cc_97 N_VSS_c_108_n N_BI_c_241_n 9.87959e-19
cc_98 N_VSS_c_119_n N_BI_c_241_n 5.43103e-19
cc_99 N_VSS_c_96_n N_BI_c_249_n 4.76944e-19
cc_100 N_VSS_c_119_n N_BI_c_249_n 6.52328e-19
cc_101 N_VSS_c_125_p N_AI_c_301_n 3.43419e-19
cc_102 N_VSS_c_97_n N_AI_c_301_n 3.48267e-19
cc_103 N_VSS_c_125_p N_AI_c_303_n 3.48267e-19
cc_104 N_VSS_c_92_n N_AI_c_303_n 0.00173332f
cc_105 N_VSS_c_97_n N_AI_c_303_n 0.00144307f
cc_106 N_VSS_c_108_n N_AI_c_303_n 0.00107717f
cc_107 N_VSS_c_97_n N_AI_c_306_n 0.0019327f
cc_108 N_VSS_c_100_n N_AI_c_306_n 0.0067288f
cc_109 N_VSS_c_97_n N_AI_c_315_n 2.82216e-19
cc_110 N_VSS_c_100_n N_AI_c_316_n 0.00177928f
cc_111 N_VSS_XI11.X0_PGD N_B_c_341_n 3.95536e-19
cc_112 N_VSS_c_108_n N_B_c_342_n 7.63393e-19
cc_113 N_VSS_c_96_n N_B_c_351_n 5.01254e-19
cc_114 N_VSS_c_125_p N_C_c_409_n 3.43419e-19
cc_115 N_VSS_c_125_p N_C_c_410_n 3.48267e-19
cc_116 N_VSS_c_97_n N_C_c_410_n 6.01757e-19
cc_117 N_A_c_187_p N_BI_XI15.X0_CG 2.06538e-19
cc_118 N_A_XI14.X0_PGD N_BI_c_252_n 9.65637e-19
cc_119 N_A_c_162_n N_BI_c_241_n 3.93183e-19
cc_120 N_A_c_179_n N_BI_c_241_n 3.15833e-19
cc_121 N_A_c_179_n N_BI_c_249_n 0.00163472f
cc_122 N_A_c_187_p N_BI_c_249_n 8.66815e-19
cc_123 N_A_c_187_p N_BI_c_257_n 4.7863e-19
cc_124 N_A_c_179_n N_BI_c_258_n 3.37713e-19
cc_125 N_A_XI14.X0_PGD N_BI_c_259_n 0.00245019f
cc_126 N_A_c_187_p N_BI_c_260_n 0.00112715f
cc_127 N_A_c_162_n N_BI_c_261_n 7.8464e-19
cc_128 N_A_XI14.X0_PGD N_AI_XI15.X0_PGD 0.0173811f
cc_129 N_A_c_179_n N_AI_XI15.X0_PGD 7.90282e-19
cc_130 N_A_c_187_p N_AI_XI15.X0_PGD 0.00103582f
cc_131 N_A_c_201_p N_AI_c_299_n 0.00196947f
cc_132 N_A_c_187_p N_AI_c_299_n 9.91291e-19
cc_133 N_A_c_203_p N_AI_c_300_n 0.00200674f
cc_134 N_A_c_161_n N_AI_c_301_n 7.16634e-19
cc_135 N_A_c_162_n N_AI_c_303_n 8.04759e-19
cc_136 N_A_c_162_n N_AI_c_306_n 0.00148587f
cc_137 N_A_XI14.X0_PGD N_B_XI14.X0_CG 9.65637e-19
cc_138 N_A_c_161_n N_B_c_341_n 0.00297252f
cc_139 N_A_c_162_n N_B_c_341_n 5.2287e-19
cc_140 N_A_c_170_n N_B_c_355_n 4.73714e-19
cc_141 N_A_c_179_n N_B_c_342_n 5.60543e-19
cc_142 N_A_c_162_n B 0.00101165f
cc_143 N_A_c_179_n B 7.63651e-19
cc_144 N_A_c_187_p N_B_c_359_n 3.89825e-19
cc_145 N_A_c_215_p N_B_c_359_n 7.82672e-19
cc_146 N_A_c_216_p N_B_c_359_n 3.42845e-19
cc_147 N_A_c_161_n N_B_c_346_n 0.00100571f
cc_148 N_A_c_179_n N_B_c_346_n 2.04384e-19
cc_149 N_A_XI14.X0_PGD N_B_c_364_n 0.00312702f
cc_150 N_A_c_216_p N_B_c_364_n 2.56268e-19
cc_151 N_A_c_162_n N_B_c_351_n 0.00214888f
cc_152 N_A_c_179_n N_B_c_351_n 0.00203212f
cc_153 N_A_c_223_p N_B_c_351_n 3.75372e-19
cc_154 N_A_c_187_p N_B_c_351_n 5.5912e-19
cc_155 N_A_c_162_n N_B_c_370_n 4.2957e-19
cc_156 N_A_c_162_n N_B_c_371_n 2.29222e-19
cc_157 N_A_c_172_n N_Z_c_427_n 3.43419e-19
cc_158 N_A_c_228_p N_Z_c_427_n 3.43419e-19
cc_159 N_A_c_223_p N_Z_c_427_n 3.48267e-19
cc_160 N_A_c_230_p N_Z_c_427_n 3.48267e-19
cc_161 N_A_c_187_p N_Z_c_427_n 7.95142e-19
cc_162 N_A_XI14.X0_PGD N_Z_c_432_n 6.68421e-19
cc_163 N_A_c_172_n N_Z_c_432_n 3.48267e-19
cc_164 N_A_c_228_p N_Z_c_432_n 3.48267e-19
cc_165 N_A_c_179_n N_Z_c_432_n 0.00126628f
cc_166 N_A_c_223_p N_Z_c_432_n 7.9714e-19
cc_167 N_A_c_230_p N_Z_c_432_n 8.16241e-19
cc_168 N_A_c_187_p N_Z_c_432_n 0.00136994f
cc_169 N_BI_XI15.X0_CG N_AI_XI15.X0_PGD 9.47088e-19
cc_170 N_BI_c_258_n N_AI_XI15.X0_PGD 0.00312702f
cc_171 N_BI_c_261_n N_AI_c_303_n 3.29431e-19
cc_172 N_BI_c_249_n N_AI_c_306_n 3.35097e-19
cc_173 N_BI_c_239_n N_B_c_341_n 9.28554e-19
cc_174 N_BI_c_249_n N_B_c_342_n 0.00169958f
cc_175 N_BI_c_249_n N_B_c_374_n 7.4385e-19
cc_176 N_BI_c_257_n N_B_c_359_n 0.00182538f
cc_177 N_BI_c_259_n N_B_c_359_n 4.99367e-19
cc_178 N_BI_c_260_n N_B_c_359_n 0.00165504f
cc_179 N_BI_c_258_n N_B_c_378_n 0.00520211f
cc_180 N_BI_c_259_n N_B_c_378_n 7.2092e-19
cc_181 N_BI_c_257_n N_B_c_364_n 4.99367e-19
cc_182 N_BI_c_258_n N_B_c_364_n 6.22265e-19
cc_183 N_BI_c_259_n N_B_c_364_n 0.00494186f
cc_184 N_BI_c_249_n N_B_c_351_n 0.00529659f
cc_185 N_BI_c_249_n N_B_c_371_n 2.67017e-19
cc_186 N_BI_c_260_n N_B_c_371_n 0.0013533f
cc_187 N_BI_c_280_p N_B_c_371_n 0.00340518f
cc_188 N_BI_c_249_n N_B_c_387_n 4.99817e-19
cc_189 N_BI_c_260_n N_B_c_387_n 9.41136e-19
cc_190 N_BI_c_283_p N_B_c_387_n 7.35033e-19
cc_191 N_BI_c_280_p N_B_c_390_n 0.00181541f
cc_192 N_BI_c_249_n N_B_c_391_n 0.00145499f
cc_193 N_BI_c_260_n N_B_c_391_n 8.66399e-19
cc_194 N_BI_c_249_n N_C_c_412_n 0.00107247f
cc_195 N_BI_c_257_n N_C_c_412_n 0.00130194f
cc_196 N_BI_c_283_p N_C_c_412_n 3.02033e-19
cc_197 N_BI_c_249_n N_Z_c_432_n 0.00190811f
cc_198 N_BI_c_257_n N_Z_c_432_n 0.00192905f
cc_199 N_BI_c_258_n N_Z_c_432_n 8.66889e-19
cc_200 N_BI_c_259_n N_Z_c_432_n 8.66889e-19
cc_201 N_BI_c_260_n N_Z_c_432_n 0.00107118f
cc_202 N_BI_c_280_p N_Z_c_432_n 0.00210701f
cc_203 N_BI_c_283_p N_Z_c_432_n 0.00100479f
cc_204 N_AI_XI15.X0_PGD N_B_c_393_n 9.65637e-19
cc_205 N_AI_c_306_n N_B_c_374_n 4.95395e-19
cc_206 N_AI_c_315_n N_B_c_374_n 3.42845e-19
cc_207 N_AI_XI15.X0_PGD N_B_c_378_n 0.00312702f
cc_208 N_AI_c_315_n N_B_c_378_n 2.56268e-19
cc_209 N_AI_c_306_n N_B_c_351_n 0.00314548f
cc_210 N_AI_c_306_n N_B_c_370_n 2.5452e-19
cc_211 N_AI_c_306_n N_B_c_371_n 2.35352e-19
cc_212 N_AI_c_306_n N_C_c_410_n 0.00152957f
cc_213 N_AI_c_306_n N_C_c_412_n 0.0018056f
cc_214 N_AI_XI15.X0_PGD N_Z_c_432_n 3.73496e-19
cc_215 N_B_c_351_n N_C_c_410_n 5.20324e-19
cc_216 N_B_c_359_n N_C_c_412_n 9.16187e-19
cc_217 N_B_c_351_n N_C_c_412_n 3.71107e-19
cc_218 N_B_c_387_n N_C_c_412_n 0.00455868f
cc_219 N_B_c_374_n N_Z_c_432_n 0.00210508f
cc_220 N_B_c_359_n N_Z_c_432_n 0.0019232f
cc_221 N_B_c_364_n N_Z_c_432_n 8.66889e-19
cc_222 N_B_c_371_n N_Z_c_432_n 4.75654e-19
cc_223 N_C_c_409_n N_Z_c_451_n 3.43419e-19
cc_224 N_C_c_422_p N_Z_c_451_n 3.43419e-19
cc_225 N_C_c_410_n N_Z_c_451_n 3.48267e-19
cc_226 N_C_c_412_n N_Z_c_451_n 3.48267e-19
cc_227 N_C_c_410_n N_Z_c_432_n 6.20216e-19
cc_228 N_C_c_412_n N_Z_c_432_n 0.00126042f
*
.ends
*
*
.subckt MAJ3_HPNW8 A B C Y VDD VSS
xgate (VDD VSS A B C Y) G4_MAJ3_N2
.ends
*
* File: G3_MIN3_T6_N2.pex.netlist
* Created: Fri Apr  1 16:54:39 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MIN3_T6_N2_VSS 2 4 6 8 10 12 27 32 37 40 42 45 53 57 60 65 70 75
+ 88 89 93 99 101 106 109 Vss
c66 107 Vss 6.43136e-19
c67 106 Vss 0.0038619f
c68 101 Vss 0.00207473f
c69 99 Vss 0.0082602f
c70 94 Vss 0.00137551f
c71 93 Vss 0.00772839f
c72 89 Vss 6.57551e-19
c73 88 Vss 0.00490261f
c74 75 Vss 0.00537019f
c75 70 Vss 7.10513e-22
c76 65 Vss 0.00231683f
c77 60 Vss 0.00177007f
c78 57 Vss 0.00552514f
c79 53 Vss 0.00488234f
c80 45 Vss 0.0850774f
c81 42 Vss 0.0849587f
c82 37 Vss 0.0679309f
c83 32 Vss 0.103906f
c84 27 Vss 0.307039f
c85 22 Vss 0.141189f
c86 10 Vss 0.134855f
c87 8 Vss 0.00171956f
c88 6 Vss 0.135276f
c89 2 Vss 0.134005f
r90 106 109 0.326018
r91 105 106 4.58464
r92 101 105 0.655813
r93 100 107 0.494161
r94 99 109 0.326018
r95 99 100 13.0037
r96 95 107 0.128424
r97 93 107 0.494161
r98 93 94 10.0862
r99 88 94 0.652036
r100 87 89 0.655813
r101 87 88 12.7536
r102 70 101 1.82344
r103 65 95 5.2515
r104 60 75 1.16709
r105 60 89 1.82344
r106 57 70 1.16709
r107 53 65 1.16709
r108 45 47 1.8672
r109 42 44 1.8672
r110 40 75 0.50025
r111 37 40 1.92555
r112 33 47 0.0685365
r113 32 34 0.652036
r114 32 33 2.8008
r115 29 47 0.5835
r116 28 42 0.0685365
r117 27 45 0.0685365
r118 27 28 10.9698
r119 24 44 0.5835
r120 23 37 0.0685365
r121 22 44 0.0685365
r122 22 23 4.7847
r123 12 57 0.185659
r124 10 34 3.8511
r125 8 53 0.185659
r126 6 29 3.8511
r127 4 53 0.185659
r128 2 24 3.8511
.ends

.subckt PM_G3_MIN3_T6_N2_VDD 2 4 6 8 10 12 27 32 42 45 53 57 60 61 63 65 69 71
+ 73 78 81 83 Vss
c76 83 Vss 0.00671487f
c77 79 Vss 7.78098e-19
c78 78 Vss 0.00468194f
c79 73 Vss 0.00129457f
c80 71 Vss 0.0122041f
c81 69 Vss 0.00238015f
c82 65 Vss 0.00185683f
c83 63 Vss 7.50392e-19
c84 62 Vss 0.0017907f
c85 61 Vss 0.007913f
c86 60 Vss 0.00707888f
c87 57 Vss 0.00500133f
c88 53 Vss 0.00483876f
c89 45 Vss 0.0849087f
c90 42 Vss 0.0854801f
c91 38 Vss 0.0711342f
c92 32 Vss 0.106714f
c93 27 Vss 0.308162f
c94 22 Vss 0.144473f
c95 12 Vss 0.13249f
c96 8 Vss 0.133305f
c97 6 Vss 0.00171956f
c98 4 Vss 0.133098f
r99 78 81 0.349767
r100 77 78 4.58464
r101 73 81 0.306046
r102 73 75 1.82344
r103 72 79 0.494161
r104 71 77 0.652036
r105 71 72 13.0037
r106 67 79 0.128424
r107 67 69 5.2515
r108 65 83 1.16709
r109 63 65 1.82344
r110 61 79 0.494161
r111 61 62 10.0862
r112 60 63 0.655813
r113 59 62 0.652036
r114 59 60 12.7536
r115 57 75 1.16709
r116 53 69 1.16709
r117 45 46 1.8672
r118 42 43 1.8672
r119 38 83 0.50025
r120 38 40 1.92555
r121 33 45 0.0685365
r122 32 34 0.652036
r123 32 33 2.8008
r124 29 45 0.5835
r125 28 43 0.0685365
r126 27 46 0.0685365
r127 27 28 10.9698
r128 24 42 0.5835
r129 23 40 0.0685365
r130 22 42 0.0685365
r131 22 23 4.7847
r132 12 34 3.8511
r133 10 57 0.185659
r134 8 29 3.8511
r135 6 53 0.185659
r136 4 24 3.8511
r137 2 53 0.185659
.ends

.subckt PM_G3_MIN3_T6_N2_Z 2 4 6 8 10 12 32 36 41 45 49 53 55 59 63 67 Vss
c60 67 Vss 3.51451e-19
c61 65 Vss 2.45386e-19
c62 63 Vss 0.00102688f
c63 59 Vss 7.58182e-19
c64 55 Vss 0.00456155f
c65 53 Vss 6.51205e-19
c66 49 Vss 6.88903e-19
c67 45 Vss 0.00781677f
c68 41 Vss 0.00689463f
c69 36 Vss 0.00387467f
c70 32 Vss 0.00319091f
c71 12 Vss 0.00171956f
c72 10 Vss 0.00171956f
r73 61 67 0.494161
r74 61 63 3.04254
r75 57 67 0.494161
r76 57 59 3.04254
r77 56 65 0.128424
r78 55 67 0.128424
r79 55 56 10.3363
r80 51 65 0.494161
r81 51 53 3.04254
r82 47 65 0.494161
r83 47 49 3.04254
r84 45 63 1.16709
r85 41 59 1.16709
r86 36 53 1.16709
r87 32 49 1.16709
r88 12 45 0.185659
r89 10 41 0.185659
r90 8 45 0.185659
r91 6 41 0.185659
r92 4 36 0.185659
r93 2 32 0.185659
.ends

.subckt PM_G3_MIN3_T6_N2_C 2 4 6 8 14 20 26 29 33 38 43 Vss
c35 43 Vss 0.00523941f
c36 38 Vss 0.00156891f
c37 33 Vss 0.00543691f
c38 29 Vss 3.56438e-22
c39 20 Vss 0.377731f
c40 14 Vss 0.380603f
r41 33 43 1.16709
r42 29 38 1.16709
r43 29 33 10.0654
r44 26 29 0.0729375
r45 20 43 0.50025
r46 14 38 0.50025
r47 6 8 10.1529
r48 6 20 3.09255
r49 2 4 10.1529
r50 2 14 3.09255
.ends

.subckt PM_G3_MIN3_T6_N2_B 2 4 6 8 17 18 26 29 35 Vss
c31 35 Vss 0.00144085f
c32 26 Vss 0.0839596f
c33 18 Vss 0.0346166f
c34 17 Vss 0.0963518f
c35 6 Vss 0.399392f
c36 2 Vss 0.447969f
r37 32 35 1.16709
r38 29 32 0.0833571
r39 24 35 0.0476429
r40 24 26 1.92555
r41 17 19 0.652036
r42 17 18 2.8008
r43 14 26 0.0685365
r44 13 18 0.652036
r45 6 8 10.1529
r46 6 19 3.8511
r47 4 14 3.8511
r48 2 4 10.1529
r49 2 13 3.8511
.ends

.subckt PM_G3_MIN3_T6_N2_A 2 4 6 8 17 29 34 38 41 46 Vss
c28 46 Vss 0.00532741f
c29 41 Vss 0.00134116f
c30 34 Vss 0.00178881f
c31 26 Vss 0.0871242f
c32 6 Vss 0.406031f
c33 2 Vss 0.376065f
r34 34 46 1.16709
r35 34 38 0.0416786
r36 29 41 1.16709
r37 29 34 5.03269
r38 24 46 0.0476429
r39 24 26 1.92555
r40 19 26 0.0685365
r41 17 41 0.50025
r42 8 19 3.8511
r43 6 8 10.1529
r44 4 17 3.09255
r45 2 4 10.1529
.ends

.subckt G3_MIN3_T6_N2  VSS VDD Z C B A
*
* A	A
* B	B
* C	C
* Z	Z
* VDD	VDD
* VSS	VSS
XI17.X0 N_Z_XI17.X0_D N_VSS_XI17.X0_PGD N_C_XI17.X0_CG N_B_XI17.X0_PGS
+ N_VDD_XI17.X0_S TIGFET_HPNW8
XI14.X0 N_Z_XI14.X0_D N_VDD_XI14.X0_PGD N_C_XI14.X0_CG N_B_XI14.X0_PGS
+ N_VSS_XI14.X0_S TIGFET_HPNW8
XI19.X0 N_Z_XI19.X0_D N_VSS_XI19.X0_PGD N_A_XI19.X0_CG N_B_XI19.X0_PGS
+ N_VDD_XI19.X0_S TIGFET_HPNW8
XI16.X0 N_Z_XI16.X0_D N_VDD_XI16.X0_PGD N_A_XI16.X0_CG N_B_XI16.X0_PGS
+ N_VSS_XI16.X0_S TIGFET_HPNW8
XI18.X0 N_Z_XI18.X0_D N_VSS_XI18.X0_PGD N_C_XI18.X0_CG N_A_XI18.X0_PGS
+ N_VDD_XI18.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_VDD_XI15.X0_PGD N_C_XI15.X0_CG N_A_XI15.X0_PGS
+ N_VSS_XI15.X0_S TIGFET_HPNW8
*
x_PM_G3_MIN3_T6_N2_VSS N_VSS_XI17.X0_PGD N_VSS_XI14.X0_S N_VSS_XI19.X0_PGD
+ N_VSS_XI16.X0_S N_VSS_XI18.X0_PGD N_VSS_XI15.X0_S N_VSS_c_19_p N_VSS_c_21_p
+ N_VSS_c_7_p N_VSS_c_13_p N_VSS_c_14_p N_VSS_c_50_p N_VSS_c_4_p N_VSS_c_22_p
+ N_VSS_c_8_p N_VSS_c_28_p N_VSS_c_6_p N_VSS_c_9_p N_VSS_c_10_p N_VSS_c_11_p
+ N_VSS_c_18_p N_VSS_c_47_p N_VSS_c_24_p N_VSS_c_66_p VSS Vss
+ PM_G3_MIN3_T6_N2_VSS
x_PM_G3_MIN3_T6_N2_VDD N_VDD_XI17.X0_S N_VDD_XI14.X0_PGD N_VDD_XI19.X0_S
+ N_VDD_XI16.X0_PGD N_VDD_XI18.X0_S N_VDD_XI15.X0_PGD N_VDD_c_70_n N_VDD_c_141_p
+ N_VDD_c_134_p N_VDD_c_133_p N_VDD_c_71_n N_VDD_c_72_n N_VDD_c_73_n
+ N_VDD_c_78_n N_VDD_c_82_n N_VDD_c_83_n N_VDD_c_85_n N_VDD_c_86_n N_VDD_c_88_n
+ N_VDD_c_123_p VDD N_VDD_c_91_n Vss PM_G3_MIN3_T6_N2_VDD
x_PM_G3_MIN3_T6_N2_Z N_Z_XI17.X0_D N_Z_XI14.X0_D N_Z_XI19.X0_D N_Z_XI16.X0_D
+ N_Z_XI18.X0_D N_Z_XI15.X0_D N_Z_c_143_n N_Z_c_144_n N_Z_c_166_n N_Z_c_146_n
+ N_Z_c_150_n N_Z_c_152_n N_Z_c_155_n N_Z_c_180_n N_Z_c_157_n Z Vss
+ PM_G3_MIN3_T6_N2_Z
x_PM_G3_MIN3_T6_N2_C N_C_XI17.X0_CG N_C_XI14.X0_CG N_C_XI18.X0_CG N_C_XI15.X0_CG
+ N_C_c_203_n N_C_c_204_n C N_C_c_210_n N_C_c_205_n N_C_c_207_n N_C_c_208_n Vss
+ PM_G3_MIN3_T6_N2_C
x_PM_G3_MIN3_T6_N2_B N_B_XI17.X0_PGS N_B_XI14.X0_PGS N_B_XI19.X0_PGS
+ N_B_XI16.X0_PGS N_B_c_242_n N_B_c_243_n N_B_c_251_n B N_B_c_253_n Vss
+ PM_G3_MIN3_T6_N2_B
x_PM_G3_MIN3_T6_N2_A N_A_XI19.X0_CG N_A_XI16.X0_CG N_A_XI18.X0_PGS
+ N_A_XI15.X0_PGS N_A_c_283_n N_A_c_270_n N_A_c_272_n A N_A_c_278_n N_A_c_279_n
+ Vss PM_G3_MIN3_T6_N2_A
cc_1 N_VSS_XI17.X0_PGD N_VDD_XI14.X0_PGD 6.38995e-19
cc_2 N_VSS_XI19.X0_PGD N_VDD_XI16.X0_PGD 6.38995e-19
cc_3 N_VSS_XI18.X0_PGD N_VDD_XI15.X0_PGD 6.25013e-19
cc_4 N_VSS_c_4_p N_VDD_c_70_n 4.60829e-19
cc_5 N_VSS_c_4_p N_VDD_c_71_n 8.28334e-19
cc_6 N_VSS_c_6_p N_VDD_c_72_n 2.52506e-19
cc_7 N_VSS_c_7_p N_VDD_c_73_n 2.61781e-19
cc_8 N_VSS_c_8_p N_VDD_c_73_n 0.00161042f
cc_9 N_VSS_c_9_p N_VDD_c_73_n 0.00119047f
cc_10 N_VSS_c_10_p N_VDD_c_73_n 0.00515748f
cc_11 N_VSS_c_11_p N_VDD_c_73_n 0.00184852f
cc_12 N_VSS_c_7_p N_VDD_c_78_n 8.70611e-19
cc_13 N_VSS_c_13_p N_VDD_c_78_n 3.72495e-19
cc_14 N_VSS_c_14_p N_VDD_c_78_n 7.57734e-19
cc_15 N_VSS_c_8_p N_VDD_c_78_n 9.95408e-19
cc_16 N_VSS_c_10_p N_VDD_c_82_n 0.00175335f
cc_17 N_VSS_c_8_p N_VDD_c_83_n 5.25611e-19
cc_18 N_VSS_c_18_p N_VDD_c_83_n 4.37902e-19
cc_19 N_VSS_c_19_p N_VDD_c_85_n 0.00120274f
cc_20 N_VSS_c_19_p N_VDD_c_86_n 8.56547e-19
cc_21 N_VSS_c_21_p N_VDD_c_86_n 8.4058e-19
cc_22 N_VSS_c_22_p N_VDD_c_88_n 2.52506e-19
cc_23 N_VSS_c_6_p N_VDD_c_88_n 3.68696e-19
cc_24 N_VSS_c_24_p N_VDD_c_88_n 0.0014668f
cc_25 N_VSS_c_9_p N_VDD_c_91_n 5.6037e-19
cc_26 N_VSS_c_9_p N_Z_c_143_n 0.00379015f
cc_27 N_VSS_c_4_p N_Z_c_144_n 3.43419e-19
cc_28 N_VSS_c_28_p N_Z_c_144_n 3.48267e-19
cc_29 N_VSS_c_4_p N_Z_c_146_n 3.43419e-19
cc_30 N_VSS_c_22_p N_Z_c_146_n 3.43419e-19
cc_31 N_VSS_c_28_p N_Z_c_146_n 3.48267e-19
cc_32 N_VSS_c_6_p N_Z_c_146_n 3.48267e-19
cc_33 N_VSS_c_8_p N_Z_c_150_n 6.97647e-19
cc_34 N_VSS_c_10_p N_Z_c_150_n 0.00155764f
cc_35 N_VSS_c_4_p N_Z_c_152_n 3.48267e-19
cc_36 N_VSS_c_28_p N_Z_c_152_n 5.03066e-19
cc_37 N_VSS_c_18_p N_Z_c_152_n 5.19985e-19
cc_38 N_VSS_c_28_p N_Z_c_155_n 9.68887e-19
cc_39 N_VSS_c_18_p N_Z_c_155_n 2.48288e-19
cc_40 N_VSS_c_4_p N_Z_c_157_n 3.48267e-19
cc_41 N_VSS_c_22_p N_Z_c_157_n 3.48267e-19
cc_42 N_VSS_c_28_p N_Z_c_157_n 4.99861e-19
cc_43 N_VSS_c_6_p N_Z_c_157_n 5.71987e-19
cc_44 N_VSS_XI17.X0_PGD N_C_c_203_n 4.30517e-19
cc_45 N_VSS_XI18.X0_PGD N_C_c_204_n 5.02359e-19
cc_46 N_VSS_c_18_p N_C_c_205_n 2.62126e-19
cc_47 N_VSS_c_47_p N_C_c_205_n 5.86314e-19
cc_48 N_VSS_XI17.X0_PGD N_C_c_207_n 4.3583e-19
cc_49 N_VSS_XI18.X0_PGD N_C_c_208_n 3.76133e-19
cc_50 N_VSS_c_50_p N_C_c_208_n 2.17009e-19
cc_51 N_VSS_XI17.X0_PGD N_B_XI17.X0_PGS 0.00109504f
cc_52 N_VSS_XI19.X0_PGD N_B_XI17.X0_PGS 2.15671e-19
cc_53 N_VSS_XI19.X0_PGD N_B_XI19.X0_PGS 0.00177732f
cc_54 N_VSS_XI18.X0_PGD N_B_XI19.X0_PGS 2.22194e-19
cc_55 N_VSS_c_50_p N_B_c_242_n 0.00177732f
cc_56 N_VSS_c_19_p N_B_c_243_n 0.00719168f
cc_57 N_VSS_c_14_p N_B_c_243_n 0.00109504f
cc_58 N_VSS_c_28_p B 2.11465e-19
cc_59 N_VSS_c_10_p B 2.74582e-19
cc_60 N_VSS_c_18_p B 3.96756e-19
cc_61 N_VSS_c_19_p N_A_XI19.X0_CG 2.63627e-19
cc_62 N_VSS_c_28_p N_A_c_270_n 3.13396e-19
cc_63 N_VSS_c_47_p N_A_c_270_n 5.88825e-19
cc_64 N_VSS_c_28_p N_A_c_272_n 0.00159318f
cc_65 N_VSS_c_47_p N_A_c_272_n 0.00984051f
cc_66 N_VSS_c_66_p N_A_c_272_n 0.00110288f
cc_67 N_VDD_c_71_n N_Z_c_143_n 3.43419e-19
cc_68 N_VDD_c_73_n N_Z_c_143_n 3.70842e-19
cc_69 N_VDD_c_78_n N_Z_c_143_n 3.4118e-19
cc_70 N_VDD_c_85_n N_Z_c_143_n 3.48267e-19
cc_71 N_VDD_c_91_n N_Z_c_144_n 0.00379015f
cc_72 N_VDD_c_71_n N_Z_c_166_n 3.43419e-19
cc_73 N_VDD_c_72_n N_Z_c_166_n 3.43419e-19
cc_74 N_VDD_c_85_n N_Z_c_166_n 3.48267e-19
cc_75 N_VDD_c_86_n N_Z_c_166_n 3.4118e-19
cc_76 N_VDD_c_88_n N_Z_c_166_n 3.72199e-19
cc_77 N_VDD_c_71_n N_Z_c_150_n 3.48267e-19
cc_78 N_VDD_c_73_n N_Z_c_150_n 0.00302769f
cc_79 N_VDD_c_78_n N_Z_c_150_n 6.28868e-19
cc_80 N_VDD_c_85_n N_Z_c_150_n 7.10279e-19
cc_81 N_VDD_c_83_n N_Z_c_152_n 5.83135e-19
cc_82 N_VDD_c_71_n N_Z_c_155_n 6.44146e-19
cc_83 N_VDD_c_78_n N_Z_c_155_n 2.8517e-19
cc_84 N_VDD_c_85_n N_Z_c_155_n 0.00109243f
cc_85 N_VDD_c_86_n N_Z_c_155_n 5.3605e-19
cc_86 N_VDD_c_71_n N_Z_c_180_n 3.48267e-19
cc_87 N_VDD_c_72_n N_Z_c_180_n 3.48267e-19
cc_88 N_VDD_c_85_n N_Z_c_180_n 7.22734e-19
cc_89 N_VDD_c_86_n N_Z_c_180_n 4.75018e-19
cc_90 N_VDD_c_88_n N_Z_c_180_n 8.5731e-19
cc_91 N_VDD_c_73_n N_C_c_210_n 2.63478e-19
cc_92 N_VDD_c_78_n N_C_c_210_n 0.00145322f
cc_93 N_VDD_c_85_n N_C_c_210_n 0.00137559f
cc_94 N_VDD_c_73_n N_C_c_205_n 2.14517e-19
cc_95 N_VDD_c_78_n N_C_c_205_n 7.60337e-19
cc_96 N_VDD_c_85_n N_C_c_205_n 0.00216983f
cc_97 N_VDD_c_86_n N_C_c_205_n 0.00534093f
cc_98 N_VDD_c_123_p N_C_c_205_n 7.91462e-19
cc_99 N_VDD_c_78_n N_C_c_207_n 7.51813e-19
cc_100 N_VDD_c_85_n N_C_c_207_n 8.66889e-19
cc_101 N_VDD_c_85_n N_C_c_208_n 2.22969e-19
cc_102 N_VDD_c_86_n N_C_c_208_n 2.63125e-19
cc_103 N_VDD_c_123_p N_C_c_208_n 4.2857e-19
cc_104 N_VDD_XI14.X0_PGD N_B_XI17.X0_PGS 0.00135245f
cc_105 N_VDD_XI16.X0_PGD N_B_XI17.X0_PGS 4.12959e-19
cc_106 N_VDD_c_70_n N_B_XI19.X0_PGS 0.00107949f
cc_107 N_VDD_c_70_n N_B_c_251_n 0.00255555f
cc_108 N_VDD_c_133_p N_B_c_251_n 4.12959e-19
cc_109 N_VDD_c_134_p N_B_c_253_n 0.00495207f
cc_110 N_VDD_c_91_n N_B_c_253_n 4.60491e-19
cc_111 N_VDD_XI16.X0_PGD N_A_XI19.X0_CG 4.83278e-19
cc_112 N_VDD_XI15.X0_PGD N_A_XI18.X0_PGS 0.00150004f
cc_113 N_VDD_c_86_n N_A_XI18.X0_PGS 2.04873e-19
cc_114 N_VDD_XI16.X0_PGD N_A_c_278_n 5.50272e-19
cc_115 N_VDD_XI15.X0_PGD N_A_c_279_n 3.23173e-19
cc_116 N_VDD_c_141_p N_A_c_279_n 0.00145458f
cc_117 N_VDD_c_133_p N_A_c_279_n 2.17009e-19
cc_118 N_Z_c_150_n N_C_c_203_n 2.87038e-19
cc_119 N_Z_c_152_n N_C_c_203_n 2.87038e-19
cc_120 N_Z_c_155_n N_C_c_203_n 6.35192e-19
cc_121 N_Z_c_180_n N_C_c_204_n 0.00103972f
cc_122 N_Z_c_155_n N_C_c_210_n 3.21572e-19
cc_123 N_Z_c_155_n N_C_c_205_n 0.00152991f
cc_124 N_Z_c_180_n N_C_c_205_n 2.21606e-19
cc_125 N_Z_c_155_n N_C_c_207_n 5.52863e-19
cc_126 N_Z_c_155_n N_B_XI17.X0_PGS 7.14549e-19
cc_127 N_Z_c_155_n N_B_XI19.X0_PGS 7.57192e-19
cc_128 N_Z_c_155_n B 4.22756e-19
cc_129 N_Z_c_155_n N_B_c_253_n 5.52863e-19
cc_130 N_Z_c_155_n N_A_XI19.X0_CG 6.53623e-19
cc_131 N_Z_c_155_n N_A_c_283_n 2.7527e-19
cc_132 N_Z_c_155_n N_A_c_270_n 3.25192e-19
cc_133 N_Z_c_155_n N_A_c_272_n 2.57254e-19
cc_134 N_Z_c_157_n N_A_c_272_n 4.03022e-19
cc_135 N_Z_c_155_n N_A_c_278_n 2.77593e-19
cc_136 N_C_c_203_n N_B_XI17.X0_PGS 0.00849032f
cc_137 N_C_c_207_n N_B_XI17.X0_PGS 3.76133e-19
cc_138 N_C_c_203_n N_B_XI19.X0_PGS 6.67601e-19
cc_139 N_C_c_204_n N_B_XI19.X0_PGS 4.29907e-19
cc_140 N_C_c_204_n N_A_XI19.X0_CG 0.00200107f
cc_141 N_C_c_204_n N_A_XI18.X0_PGS 0.00801113f
cc_142 N_C_c_205_n N_A_c_272_n 0.00154898f
cc_143 N_B_XI17.X0_PGS N_A_XI19.X0_CG 8.40291e-19
cc_144 N_B_XI19.X0_PGS N_A_XI19.X0_CG 0.00774979f
cc_145 B N_A_c_270_n 3.39698e-19
cc_146 N_B_c_253_n N_A_c_270_n 3.48267e-19
cc_147 B N_A_c_278_n 3.48267e-19
cc_148 N_B_c_253_n N_A_c_278_n 5.15124e-19
*
.ends
*
*
.subckt MIN3_HPNW8 A B C Y VDD VSS
xgate (VSS VDD Y C B A) G3_MIN3_T6_N2
.ends
*
* File: G4_MUX2_N2.pex.netlist
* Created: Tue Mar 15 11:14:18 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MUX2_N2_VDD 2 4 6 8 10 12 14 16 18 20 38 49 51 58 64 72 77 81 84
+ 85 89 93 95 96 99 101 105 107 111 113 115 120 122 124 125 126 127 128 134 139
+ 148 Vss
c133 148 Vss 0.00699273f
c134 139 Vss 0.00445774f
c135 134 Vss 0.00494975f
c136 128 Vss 4.52364e-19
c137 127 Vss 2.39889e-19
c138 126 Vss 4.2334e-19
c139 125 Vss 2.39889e-19
c140 122 Vss 0.00207203f
c141 120 Vss 0.00831709f
c142 115 Vss 0.00192f
c143 113 Vss 0.00621353f
c144 111 Vss 7.23227e-19
c145 107 Vss 0.00783849f
c146 105 Vss 0.0013925f
c147 101 Vss 0.00172494f
c148 99 Vss 3.98903e-19
c149 96 Vss 6.1175e-19
c150 95 Vss 0.00348383f
c151 93 Vss 0.00103115f
c152 89 Vss 0.0016395f
c153 86 Vss 0.00175544f
c154 85 Vss 0.00656595f
c155 84 Vss 0.0047574f
c156 81 Vss 0.00425172f
c157 77 Vss 0.00710807f
c158 72 Vss 0.00394783f
c159 64 Vss 9.76046e-20
c160 59 Vss 0.0805856f
c161 58 Vss 0.104002f
c162 51 Vss 1.36639e-19
c163 49 Vss 0.035607f
c164 48 Vss 0.101298f
c165 39 Vss 0.0367217f
c166 38 Vss 0.101451f
c167 18 Vss 0.134291f
c168 16 Vss 0.00143442f
c169 14 Vss 0.136641f
c170 10 Vss 0.134979f
c171 8 Vss 0.134694f
c172 6 Vss 0.136393f
c173 4 Vss 0.134706f
r174 121 128 0.551426
r175 121 122 4.58464
r176 120 128 0.551426
r177 119 120 15.5878
r178 115 128 0.0828784
r179 115 117 1.82344
r180 114 127 0.494161
r181 113 119 0.652036
r182 113 114 10.1279
r183 111 148 1.16709
r184 109 127 0.128424
r185 109 111 2.16729
r186 108 126 0.494161
r187 107 122 0.652036
r188 107 108 13.0037
r189 103 126 0.128424
r190 103 105 5.2515
r191 102 125 0.494161
r192 101 127 0.494161
r193 101 102 4.58464
r194 99 139 1.16709
r195 97 125 0.128424
r196 97 99 2.16729
r197 95 126 0.494161
r198 95 96 7.46046
r199 93 134 1.16709
r200 91 96 0.652036
r201 91 93 2.16729
r202 87 124 0.306046
r203 87 89 1.82344
r204 85 125 0.494161
r205 85 86 10.1279
r206 84 124 0.349767
r207 83 86 0.652036
r208 83 84 4.58464
r209 81 117 1.16709
r210 77 105 1.16709
r211 72 89 1.16709
r212 64 148 0.0476429
r213 64 66 1.92555
r214 59 66 0.5835
r215 58 60 0.652036
r216 58 59 2.8008
r217 55 66 0.0685365
r218 51 139 0.0476429
r219 49 51 1.45875
r220 48 52 0.652036
r221 48 51 1.45875
r222 45 49 0.652036
r223 41 134 0.0476429
r224 39 41 1.45875
r225 38 42 0.652036
r226 38 41 1.45875
r227 35 39 0.652036
r228 20 81 0.185659
r229 18 60 3.8511
r230 16 77 0.185659
r231 14 55 3.8511
r232 12 77 0.185659
r233 10 52 3.8511
r234 8 45 3.8511
r235 6 35 3.8511
r236 4 42 3.8511
r237 2 72 0.185659
.ends

.subckt PM_G4_MUX2_N2_VSS 2 4 6 8 10 12 14 16 18 20 38 39 41 48 49 59 72 77 81
+ 84 89 94 99 104 109 118 123 132 141 142 146 152 153 158 164 170 172 177 179
+ 181 182 183 184 185 Vss
c128 185 Vss 4.28045e-19
c129 184 Vss 3.62111e-19
c130 183 Vss 3.88979e-19
c131 182 Vss 3.21876e-19
c132 179 Vss 0.00491274f
c133 177 Vss 0.00148831f
c134 172 Vss 0.00130997f
c135 170 Vss 0.0025874f
c136 164 Vss 0.00591751f
c137 158 Vss 0.00396568f
c138 153 Vss 5.94991e-19
c139 152 Vss 0.00255814f
c140 146 Vss 0.00513861f
c141 142 Vss 0.00102564f
c142 141 Vss 0.00403723f
c143 132 Vss 0.00811196f
c144 123 Vss 0.00369111f
c145 118 Vss 0.00399678f
c146 109 Vss 4.35064e-19
c147 104 Vss 0.00132832f
c148 99 Vss 0.00135757f
c149 94 Vss 4.3806e-19
c150 89 Vss 9.57033e-19
c151 84 Vss 0.00151444f
c152 81 Vss 0.00400382f
c153 77 Vss 0.00617013f
c154 72 Vss 0.00549529f
c155 65 Vss 0.0783825f
c156 59 Vss 0.0350566f
c157 58 Vss 0.0688416f
c158 49 Vss 0.0347733f
c159 48 Vss 0.100344f
c160 41 Vss 9.8832e-20
c161 39 Vss 0.0350852f
c162 38 Vss 0.0994129f
c163 20 Vss 0.135394f
c164 16 Vss 0.134482f
c165 14 Vss 0.00143442f
c166 12 Vss 0.134697f
c167 10 Vss 0.135146f
c168 4 Vss 0.134814f
c169 2 Vss 0.13402f
r170 178 185 0.551426
r171 178 179 15.5878
r172 177 185 0.551426
r173 176 177 4.58464
r174 172 185 0.0828784
r175 171 184 0.494161
r176 170 179 0.652036
r177 170 171 4.41793
r178 166 184 0.128424
r179 165 183 0.494161
r180 164 176 0.652036
r181 164 165 13.0037
r182 160 183 0.128424
r183 159 182 0.494161
r184 158 184 0.494161
r185 158 159 10.2946
r186 154 182 0.128424
r187 152 183 0.494161
r188 152 153 7.46046
r189 148 153 0.652036
r190 147 181 0.326018
r191 146 182 0.494161
r192 146 147 10.1279
r193 141 181 0.326018
r194 140 142 0.655813
r195 140 141 4.58464
r196 109 172 1.82344
r197 104 132 1.16709
r198 104 166 2.16729
r199 99 160 5.2515
r200 94 123 1.16709
r201 94 154 2.16729
r202 89 118 1.16709
r203 89 148 2.16729
r204 84 142 1.82344
r205 81 109 1.16709
r206 77 99 1.16709
r207 72 84 1.16709
r208 65 132 0.0476429
r209 63 65 1.8672
r210 60 63 0.0685365
r211 58 63 0.5835
r212 58 59 2.8008
r213 55 59 0.652036
r214 51 123 0.0476429
r215 49 51 1.45875
r216 48 52 0.652036
r217 48 51 1.45875
r218 45 49 0.652036
r219 41 118 0.0476429
r220 39 41 1.45875
r221 38 42 0.652036
r222 38 41 1.45875
r223 35 39 0.652036
r224 20 60 3.8511
r225 18 81 0.185659
r226 16 55 3.8511
r227 14 77 0.185659
r228 12 52 3.8511
r229 10 45 3.8511
r230 8 77 0.185659
r231 6 72 0.185659
r232 4 35 3.8511
r233 2 42 3.8511
.ends

.subckt PM_G4_MUX2_N2_ZI 2 4 6 8 10 12 27 28 43 47 50 55 60 65 81 82 91 Vss
c67 82 Vss 9.49146e-19
c68 81 Vss 0.00328207f
c69 65 Vss 0.00492924f
c70 60 Vss 0.00114673f
c71 55 Vss 0.00119934f
c72 50 Vss 0.00186152f
c73 47 Vss 0.00662602f
c74 43 Vss 0.00662602f
c75 28 Vss 0.204565f
c76 27 Vss 9.8832e-20
c77 23 Vss 0.0247918f
c78 12 Vss 0.00143442f
c79 10 Vss 0.00143442f
c80 4 Vss 0.134965f
c81 2 Vss 0.126125f
r82 87 91 0.494161
r83 83 91 0.494161
r84 81 91 0.128424
r85 81 82 13.2121
r86 77 82 0.652036
r87 60 87 4.58464
r88 55 83 5.2515
r89 50 65 1.16709
r90 50 77 2.16729
r91 47 60 1.16709
r92 43 55 1.16709
r93 31 65 0.0476429
r94 29 31 0.326018
r95 29 31 0.1167
r96 28 32 0.652036
r97 28 31 6.7686
r98 27 65 0.357321
r99 23 31 0.326018
r100 23 27 0.40845
r101 12 47 0.185659
r102 10 43 0.185659
r103 8 47 0.185659
r104 6 43 0.185659
r105 4 32 3.8511
r106 2 27 3.44265
.ends

.subckt PM_G4_MUX2_N2_Z 2 4 13 16 19 Vss
c13 16 Vss 2.38782e-19
c14 13 Vss 0.00448964f
c15 4 Vss 0.00143442f
r16 16 19 0.0416786
r17 13 16 1.16709
r18 4 13 0.185659
r19 2 13 0.185659
.ends

.subckt PM_G4_MUX2_N2_SELI 2 4 6 8 18 21 29 33 36 38 43 44 52 57 71 76 77 Vss
c77 77 Vss 8.68628e-19
c78 76 Vss 1.71087e-19
c79 71 Vss 0.00181943f
c80 57 Vss 0.00285848f
c81 52 Vss 0.00302696f
c82 44 Vss 0.00257468f
c83 43 Vss 7.72677e-19
c84 38 Vss 0.00166363f
c85 36 Vss 3.84679e-19
c86 33 Vss 0.00302237f
c87 29 Vss 0.00550884f
c88 21 Vss 0.112078f
c89 18 Vss 1.01432e-19
c90 6 Vss 0.112115f
c91 4 Vss 0.00143442f
r92 76 77 0.655813
r93 75 76 3.501
r94 71 75 0.655813
r95 43 52 1.16709
r96 43 71 2.00578
r97 43 44 0.513084
r98 38 57 1.16709
r99 38 77 2.00578
r100 36 44 7.46046
r101 31 36 0.652036
r102 31 33 7.002
r103 29 33 1.16709
r104 21 57 0.50025
r105 18 52 0.50025
r106 8 21 3.09255
r107 6 18 3.09255
r108 4 29 0.185659
r109 2 29 0.185659
.ends

.subckt PM_G4_MUX2_N2_SEL 2 4 6 8 16 17 22 26 33 36 40 41 44 45 47 49 56 57 59
+ 64 69 Vss
c70 69 Vss 0.00270368f
c71 64 Vss 0.00315728f
c72 59 Vss 0.00270998f
c73 57 Vss 3.45787e-19
c74 56 Vss 0.00198364f
c75 49 Vss 3.06667e-19
c76 47 Vss 0.00132431f
c77 45 Vss 4.54881e-19
c78 44 Vss 0.00192809f
c79 41 Vss 0.00173298f
c80 36 Vss 9.81095e-20
c81 33 Vss 1.05421e-19
c82 26 Vss 0.112078f
c83 22 Vss 0.125771f
c84 20 Vss 0.0247918f
c85 17 Vss 0.0358516f
c86 16 Vss 0.176172f
c87 8 Vss 0.112078f
c88 2 Vss 0.139232f
r89 55 64 1.16709
r90 55 57 0.4602
r91 55 56 0.52504
r92 52 59 1.16709
r93 49 52 0.5835
r94 47 69 1.16709
r95 45 47 2.00578
r96 43 45 0.655813
r97 43 44 3.501
r98 41 44 0.655813
r99 41 57 1.49522
r100 40 56 3.04254
r101 38 49 0.0685365
r102 38 40 1.54211
r103 36 59 0.0476429
r104 33 69 0.50025
r105 26 64 0.50025
r106 22 59 0.357321
r107 20 36 0.326018
r108 20 22 0.40845
r109 17 36 6.7686
r110 16 36 0.326018
r111 16 36 0.1167
r112 13 17 0.652036
r113 8 33 3.09255
r114 6 26 3.09255
r115 4 22 3.44265
r116 2 13 3.8511
.ends

.subckt PM_G4_MUX2_N2_B 2 4 14 20 23 Vss
c30 23 Vss 0.00425113f
c31 20 Vss 3.02878e-19
c32 14 Vss 0.0853035f
c33 2 Vss 0.547212f
r34 17 23 1.16709
r35 17 20 0.0729375
r36 14 23 0.0476429
r37 11 14 1.92555
r38 7 11 0.0685365
r39 4 7 3.8511
r40 2 4 15.4044
.ends

.subckt PM_G4_MUX2_N2_A 2 4 12 14 17 23 Vss
c24 23 Vss 0.00254505f
c25 17 Vss 3.13475e-19
c26 14 Vss 0.0661045f
c27 12 Vss 1.05421e-19
c28 2 Vss 0.578847f
r29 20 23 1.16709
r30 17 20 0.0833571
r31 12 23 0.3335
r32 12 14 1.57545
r33 7 14 0.0685365
r34 2 4 15.4044
r35 2 7 4.60965
.ends

.subckt G4_MUX2_N2  VDD VSS Z SEL B A
*
* A	A
* B	B
* SEL	SEL
* Z	Z
* VSS	VSS
* VDD	VDD
XI5.X0 N_Z_XI5.X0_D N_VSS_XI5.X0_PGD N_ZI_XI5.X0_CG N_VSS_XI5.X0_PGS
+ N_VDD_XI5.X0_S TIGFET_HPNW8
XI6.X0 N_SELI_XI6.X0_D N_VDD_XI6.X0_PGD N_SEL_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VDD_XI4.X0_PGD N_ZI_XI4.X0_CG N_VDD_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW8
XI7.X0 N_SELI_XI7.X0_D N_VSS_XI7.X0_PGD N_SEL_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW8
XI11.X0 N_ZI_XI11.X0_D N_VDD_XI11.X0_PGD N_SELI_XI11.X0_CG N_B_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW8
XI9.X0 N_ZI_XI9.X0_D N_VSS_XI9.X0_PGD N_SEL_XI9.X0_CG N_B_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW8
XI10.X0 N_ZI_XI10.X0_D N_VDD_XI10.X0_PGD N_SEL_XI10.X0_CG N_A_XI10.X0_PGS
+ N_VSS_XI10.X0_S TIGFET_HPNW8
XI8.X0 N_ZI_XI8.X0_D N_VSS_XI8.X0_PGD N_SELI_XI8.X0_CG N_A_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW8
*
x_PM_G4_MUX2_N2_VDD N_VDD_XI5.X0_S N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS
+ N_VDD_XI4.X0_PGD N_VDD_XI4.X0_PGS N_VDD_XI7.X0_S N_VDD_XI11.X0_PGD
+ N_VDD_XI9.X0_S N_VDD_XI10.X0_PGD N_VDD_XI8.X0_S N_VDD_c_12_p N_VDD_c_8_p
+ N_VDD_c_115_p N_VDD_c_121_p N_VDD_c_91_p N_VDD_c_85_p N_VDD_c_15_p
+ N_VDD_c_72_p N_VDD_c_10_p N_VDD_c_9_p N_VDD_c_17_p N_VDD_c_22_p N_VDD_c_13_p
+ N_VDD_c_47_p N_VDD_c_20_p N_VDD_c_27_p N_VDD_c_5_p N_VDD_c_14_p N_VDD_c_28_p
+ N_VDD_c_16_p N_VDD_c_59_p N_VDD_c_29_p N_VDD_c_32_p VDD N_VDD_c_50_p
+ N_VDD_c_54_p N_VDD_c_57_p N_VDD_c_64_p N_VDD_c_25_p N_VDD_c_21_p N_VDD_c_100_p
+ Vss PM_G4_MUX2_N2_VDD
x_PM_G4_MUX2_N2_VSS N_VSS_XI5.X0_PGD N_VSS_XI5.X0_PGS N_VSS_XI6.X0_S
+ N_VSS_XI4.X0_S N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS N_VSS_XI11.X0_S
+ N_VSS_XI9.X0_PGD N_VSS_XI10.X0_S N_VSS_XI8.X0_PGD N_VSS_c_141_n N_VSS_c_143_n
+ N_VSS_c_202_p N_VSS_c_252_p N_VSS_c_145_n N_VSS_c_147_n N_VSS_c_227_p
+ N_VSS_c_148_n N_VSS_c_149_n N_VSS_c_150_n N_VSS_c_151_n N_VSS_c_155_n
+ N_VSS_c_159_n N_VSS_c_163_n N_VSS_c_166_n N_VSS_c_168_n N_VSS_c_171_n
+ N_VSS_c_175_n N_VSS_c_177_n N_VSS_c_178_n N_VSS_c_179_n N_VSS_c_181_n
+ N_VSS_c_184_n N_VSS_c_185_n N_VSS_c_188_n N_VSS_c_191_n N_VSS_c_192_n
+ N_VSS_c_193_n N_VSS_c_194_n VSS N_VSS_c_198_n N_VSS_c_199_n N_VSS_c_200_n
+ N_VSS_c_201_n Vss PM_G4_MUX2_N2_VSS
x_PM_G4_MUX2_N2_ZI N_ZI_XI5.X0_CG N_ZI_XI4.X0_CG N_ZI_XI11.X0_D N_ZI_XI9.X0_D
+ N_ZI_XI10.X0_D N_ZI_XI8.X0_D N_ZI_c_278_n N_ZI_c_262_n N_ZI_c_263_n
+ N_ZI_c_264_n N_ZI_c_283_n N_ZI_c_269_n N_ZI_c_271_n N_ZI_c_276_n N_ZI_c_277_n
+ N_ZI_c_298_n N_ZI_c_314_p Vss PM_G4_MUX2_N2_ZI
x_PM_G4_MUX2_N2_Z N_Z_XI5.X0_D N_Z_XI4.X0_D N_Z_c_329_n N_Z_c_332_n Z Vss
+ PM_G4_MUX2_N2_Z
x_PM_G4_MUX2_N2_SELI N_SELI_XI6.X0_D N_SELI_XI7.X0_D N_SELI_XI11.X0_CG
+ N_SELI_XI8.X0_CG N_SELI_c_342_n N_SELI_c_417_p N_SELI_c_343_n N_SELI_c_346_n
+ N_SELI_c_374_n N_SELI_c_349_n N_SELI_c_350_n N_SELI_c_352_n N_SELI_c_356_n
+ N_SELI_c_368_n N_SELI_c_370_n N_SELI_c_384_n N_SELI_c_387_n Vss
+ PM_G4_MUX2_N2_SELI
x_PM_G4_MUX2_N2_SEL N_SEL_XI6.X0_CG N_SEL_XI7.X0_CG N_SEL_XI9.X0_CG
+ N_SEL_XI10.X0_CG N_SEL_c_419_n N_SEL_c_439_n N_SEL_c_473_p N_SEL_c_474_p
+ N_SEL_c_484_p N_SEL_c_430_n SEL N_SEL_c_420_n N_SEL_c_421_n N_SEL_c_446_n
+ N_SEL_c_422_n N_SEL_c_433_n N_SEL_c_425_n N_SEL_c_462_n N_SEL_c_427_n
+ N_SEL_c_465_n N_SEL_c_428_n Vss PM_G4_MUX2_N2_SEL
x_PM_G4_MUX2_N2_B N_B_XI11.X0_PGS N_B_XI9.X0_PGS N_B_c_495_n B N_B_c_491_n Vss
+ PM_G4_MUX2_N2_B
x_PM_G4_MUX2_N2_A N_A_XI10.X0_PGS N_A_XI8.X0_PGS N_A_c_537_n N_A_c_521_n A
+ N_A_c_527_n Vss PM_G4_MUX2_N2_A
cc_1 N_VDD_XI4.X0_PGD N_VSS_XI5.X0_PGD 0.00201121f
cc_2 N_VDD_XI6.X0_PGS N_VSS_XI5.X0_PGS 2.37403e-19
cc_3 N_VDD_XI6.X0_PGD N_VSS_XI7.X0_PGD 0.00195824f
cc_4 N_VDD_XI4.X0_PGS N_VSS_XI7.X0_PGS 2.20829e-19
cc_5 N_VDD_c_5_p N_VSS_XI7.X0_PGS 2.10824e-19
cc_6 N_VDD_XI11.X0_PGD N_VSS_XI9.X0_PGD 2.24862e-19
cc_7 N_VDD_XI10.X0_PGD N_VSS_XI8.X0_PGD 2.24862e-19
cc_8 N_VDD_c_8_p N_VSS_c_141_n 0.00201121f
cc_9 N_VDD_c_9_p N_VSS_c_141_n 3.9313e-19
cc_10 N_VDD_c_10_p N_VSS_c_143_n 3.05236e-19
cc_11 N_VDD_c_9_p N_VSS_c_143_n 4.1253e-19
cc_12 N_VDD_c_12_p N_VSS_c_145_n 0.00195824f
cc_13 N_VDD_c_13_p N_VSS_c_145_n 3.03215e-19
cc_14 N_VDD_c_14_p N_VSS_c_147_n 8.80211e-19
cc_15 N_VDD_c_15_p N_VSS_c_148_n 3.1188e-19
cc_16 N_VDD_c_16_p N_VSS_c_149_n 3.4118e-19
cc_17 N_VDD_c_17_p N_VSS_c_150_n 5.69928e-19
cc_18 N_VDD_c_10_p N_VSS_c_151_n 8.67538e-19
cc_19 N_VDD_c_9_p N_VSS_c_151_n 0.00161703f
cc_20 N_VDD_c_20_p N_VSS_c_151_n 8.83788e-19
cc_21 N_VDD_c_21_p N_VSS_c_151_n 3.48267e-19
cc_22 N_VDD_c_22_p N_VSS_c_155_n 8.50587e-19
cc_23 N_VDD_c_13_p N_VSS_c_155_n 0.00161703f
cc_24 N_VDD_c_5_p N_VSS_c_155_n 0.00180638f
cc_25 N_VDD_c_25_p N_VSS_c_155_n 3.48267e-19
cc_26 N_VDD_c_20_p N_VSS_c_159_n 3.92901e-19
cc_27 N_VDD_c_27_p N_VSS_c_159_n 4.34701e-19
cc_28 N_VDD_c_28_p N_VSS_c_159_n 7.06793e-19
cc_29 N_VDD_c_29_p N_VSS_c_159_n 3.47458e-19
cc_30 N_VDD_c_5_p N_VSS_c_163_n 2.93442e-19
cc_31 N_VDD_c_14_p N_VSS_c_163_n 0.00161703f
cc_32 N_VDD_c_32_p N_VSS_c_163_n 4.28751e-19
cc_33 N_VDD_c_16_p N_VSS_c_166_n 4.19648e-19
cc_34 N_VDD_c_29_p N_VSS_c_166_n 0.00187494f
cc_35 N_VDD_c_10_p N_VSS_c_168_n 3.66936e-19
cc_36 N_VDD_c_9_p N_VSS_c_168_n 2.26455e-19
cc_37 N_VDD_c_21_p N_VSS_c_168_n 6.489e-19
cc_38 N_VDD_c_22_p N_VSS_c_171_n 3.82294e-19
cc_39 N_VDD_c_13_p N_VSS_c_171_n 2.26455e-19
cc_40 N_VDD_c_5_p N_VSS_c_171_n 9.55349e-19
cc_41 N_VDD_c_25_p N_VSS_c_171_n 6.46219e-19
cc_42 N_VDD_c_14_p N_VSS_c_175_n 2.26455e-19
cc_43 N_VDD_c_32_p N_VSS_c_175_n 3.63088e-19
cc_44 N_VDD_c_22_p N_VSS_c_177_n 3.85245e-19
cc_45 N_VDD_c_10_p N_VSS_c_178_n 4.00013e-19
cc_46 N_VDD_c_13_p N_VSS_c_179_n 0.00408997f
cc_47 N_VDD_c_47_p N_VSS_c_179_n 0.00164958f
cc_48 N_VDD_c_9_p N_VSS_c_181_n 0.0040756f
cc_49 N_VDD_c_27_p N_VSS_c_181_n 0.00132969f
cc_50 N_VDD_c_50_p N_VSS_c_181_n 0.00102696f
cc_51 N_VDD_c_9_p N_VSS_c_184_n 0.00176255f
cc_52 N_VDD_c_13_p N_VSS_c_185_n 0.00134925f
cc_53 N_VDD_c_14_p N_VSS_c_185_n 0.0059995f
cc_54 N_VDD_c_54_p N_VSS_c_185_n 0.00115121f
cc_55 N_VDD_c_27_p N_VSS_c_188_n 0.00132969f
cc_56 N_VDD_c_16_p N_VSS_c_188_n 0.00814611f
cc_57 N_VDD_c_57_p N_VSS_c_188_n 9.97418e-19
cc_58 N_VDD_c_14_p N_VSS_c_191_n 0.00456934f
cc_59 N_VDD_c_59_p N_VSS_c_192_n 4.54377e-19
cc_60 N_VDD_c_29_p N_VSS_c_193_n 0.00335336f
cc_61 N_VDD_c_5_p N_VSS_c_194_n 3.22916e-19
cc_62 N_VDD_c_29_p N_VSS_c_194_n 0.00738754f
cc_63 N_VDD_c_32_p N_VSS_c_194_n 0.00291237f
cc_64 N_VDD_c_64_p N_VSS_c_194_n 0.0010706f
cc_65 N_VDD_c_13_p N_VSS_c_198_n 7.23159e-19
cc_66 N_VDD_c_27_p N_VSS_c_199_n 0.00107375f
cc_67 N_VDD_c_14_p N_VSS_c_200_n 7.61747e-19
cc_68 N_VDD_c_29_p N_VSS_c_201_n 9.16632e-19
cc_69 N_VDD_XI4.X0_PGD N_ZI_c_262_n 3.93784e-19
cc_70 N_VDD_c_16_p N_ZI_c_263_n 3.4118e-19
cc_71 N_VDD_c_15_p N_ZI_c_264_n 3.43419e-19
cc_72 N_VDD_c_72_p N_ZI_c_264_n 3.43419e-19
cc_73 N_VDD_c_5_p N_ZI_c_264_n 3.48267e-19
cc_74 N_VDD_c_14_p N_ZI_c_264_n 3.4118e-19
cc_75 N_VDD_c_59_p N_ZI_c_264_n 3.72199e-19
cc_76 N_VDD_c_16_p N_ZI_c_269_n 3.98099e-19
cc_77 N_VDD_c_29_p N_ZI_c_269_n 7.67329e-19
cc_78 N_VDD_c_15_p N_ZI_c_271_n 3.48267e-19
cc_79 N_VDD_c_72_p N_ZI_c_271_n 3.48267e-19
cc_80 N_VDD_c_5_p N_ZI_c_271_n 4.99861e-19
cc_81 N_VDD_c_14_p N_ZI_c_271_n 3.98099e-19
cc_82 N_VDD_c_59_p N_ZI_c_271_n 5.226e-19
cc_83 N_VDD_c_25_p N_ZI_c_276_n 3.30805e-19
cc_84 N_VDD_c_13_p N_ZI_c_277_n 3.38227e-19
cc_85 N_VDD_c_85_p N_Z_c_329_n 3.43419e-19
cc_86 N_VDD_c_9_p N_Z_c_329_n 3.4118e-19
cc_87 N_VDD_c_17_p N_Z_c_329_n 3.72199e-19
cc_88 N_VDD_c_85_p N_Z_c_332_n 3.48267e-19
cc_89 N_VDD_c_9_p N_Z_c_332_n 4.58391e-19
cc_90 N_VDD_c_17_p N_Z_c_332_n 7.4527e-19
cc_91 N_VDD_c_91_p N_SELI_c_342_n 8.8401e-19
cc_92 N_VDD_c_15_p N_SELI_c_343_n 3.43419e-19
cc_93 N_VDD_c_13_p N_SELI_c_343_n 3.4118e-19
cc_94 N_VDD_c_5_p N_SELI_c_343_n 3.48267e-19
cc_95 N_VDD_c_15_p N_SELI_c_346_n 3.48267e-19
cc_96 N_VDD_c_13_p N_SELI_c_346_n 4.79144e-19
cc_97 N_VDD_c_5_p N_SELI_c_346_n 6.94315e-19
cc_98 N_VDD_c_29_p N_SELI_c_349_n 4.73641e-19
cc_99 N_VDD_c_28_p N_SELI_c_350_n 3.11429e-19
cc_100 N_VDD_c_100_p N_SELI_c_350_n 3.26631e-19
cc_101 N_VDD_XI4.X0_PGD N_SELI_c_352_n 2.33421e-19
cc_102 N_VDD_c_20_p N_SELI_c_352_n 4.24036e-19
cc_103 N_VDD_c_27_p N_SELI_c_352_n 2.6015e-19
cc_104 N_VDD_c_21_p N_SELI_c_352_n 2.91146e-19
cc_105 N_VDD_c_28_p N_SELI_c_356_n 3.43988e-19
cc_106 N_VDD_c_100_p N_SELI_c_356_n 2.68747e-19
cc_107 N_VDD_XI6.X0_PGD N_SEL_c_419_n 4.07423e-19
cc_108 N_VDD_c_14_p N_SEL_c_420_n 4.4769e-19
cc_109 N_VDD_c_29_p N_SEL_c_421_n 5.4414e-19
cc_110 N_VDD_c_14_p N_SEL_c_422_n 2.04009e-19
cc_111 N_VDD_c_16_p N_SEL_c_422_n 4.56389e-19
cc_112 N_VDD_c_29_p N_SEL_c_422_n 5.05119e-19
cc_113 N_VDD_c_15_p N_SEL_c_425_n 6.34806e-19
cc_114 N_VDD_c_5_p N_SEL_c_425_n 0.0010174f
cc_115 N_VDD_c_115_p N_SEL_c_427_n 4.97707e-19
cc_116 N_VDD_c_29_p N_SEL_c_428_n 3.66936e-19
cc_117 N_VDD_c_5_p B 0.00142218f
cc_118 N_VDD_c_14_p B 0.00141439f
cc_119 N_VDD_c_5_p N_B_c_491_n 9.67317e-19
cc_120 N_VDD_c_14_p N_B_c_491_n 0.00120343f
cc_121 N_VDD_c_121_p N_A_XI10.X0_PGS 0.00270087f
cc_122 N_VDD_c_29_p N_A_XI10.X0_PGS 0.00113883f
cc_123 N_VDD_c_16_p N_A_c_521_n 3.83429e-19
cc_124 N_VDD_c_29_p N_A_c_521_n 4.45055e-19
cc_125 N_VDD_c_28_p A 5.39847e-19
cc_126 N_VDD_c_16_p A 0.00141439f
cc_127 N_VDD_c_29_p A 4.93619e-19
cc_128 N_VDD_c_100_p A 3.48267e-19
cc_129 N_VDD_XI10.X0_PGD N_A_c_527_n 3.23173e-19
cc_130 N_VDD_c_28_p N_A_c_527_n 4.07426e-19
cc_131 N_VDD_c_16_p N_A_c_527_n 0.00124433f
cc_132 N_VDD_c_29_p N_A_c_527_n 3.66936e-19
cc_133 N_VDD_c_100_p N_A_c_527_n 6.47766e-19
cc_134 N_VSS_c_202_p N_ZI_c_278_n 9.69352e-19
cc_135 N_VSS_XI5.X0_PGD N_ZI_c_262_n 4.04227e-19
cc_136 N_VSS_c_148_n N_ZI_c_263_n 3.43419e-19
cc_137 N_VSS_c_149_n N_ZI_c_263_n 3.43419e-19
cc_138 N_VSS_c_166_n N_ZI_c_263_n 3.48267e-19
cc_139 N_VSS_c_151_n N_ZI_c_283_n 8.31001e-19
cc_140 N_VSS_c_168_n N_ZI_c_283_n 3.27324e-19
cc_141 N_VSS_c_148_n N_ZI_c_269_n 3.48267e-19
cc_142 N_VSS_c_149_n N_ZI_c_269_n 3.48267e-19
cc_143 N_VSS_c_159_n N_ZI_c_269_n 0.00100597f
cc_144 N_VSS_c_166_n N_ZI_c_269_n 4.40384e-19
cc_145 N_VSS_c_188_n N_ZI_c_269_n 4.67196e-19
cc_146 N_VSS_c_192_n N_ZI_c_269_n 6.1924e-19
cc_147 N_VSS_c_194_n N_ZI_c_269_n 0.0017026f
cc_148 N_VSS_c_185_n N_ZI_c_271_n 4.67196e-19
cc_149 N_VSS_c_168_n N_ZI_c_276_n 2.68747e-19
cc_150 N_VSS_c_155_n N_ZI_c_277_n 3.44104e-19
cc_151 N_VSS_c_159_n N_ZI_c_277_n 5.20154e-19
cc_152 N_VSS_c_181_n N_ZI_c_277_n 8.7206e-19
cc_153 N_VSS_c_185_n N_ZI_c_277_n 0.0012589f
cc_154 N_VSS_c_179_n N_ZI_c_298_n 9.87505e-19
cc_155 N_VSS_c_148_n N_Z_c_329_n 3.43419e-19
cc_156 N_VSS_c_159_n N_Z_c_329_n 3.48267e-19
cc_157 N_VSS_c_148_n N_Z_c_332_n 3.48267e-19
cc_158 N_VSS_c_159_n N_Z_c_332_n 7.85754e-19
cc_159 N_VSS_c_227_p N_SELI_c_343_n 3.43419e-19
cc_160 N_VSS_c_150_n N_SELI_c_343_n 3.48267e-19
cc_161 N_VSS_c_227_p N_SELI_c_346_n 3.48267e-19
cc_162 N_VSS_c_150_n N_SELI_c_346_n 5.71987e-19
cc_163 N_VSS_c_163_n N_SELI_c_349_n 7.9573e-19
cc_164 N_VSS_c_175_n N_SELI_c_349_n 3.2351e-19
cc_165 N_VSS_c_188_n N_SELI_c_349_n 4.51137e-19
cc_166 N_VSS_c_194_n N_SELI_c_349_n 6.69121e-19
cc_167 N_VSS_c_159_n N_SELI_c_352_n 0.00105826f
cc_168 N_VSS_c_181_n N_SELI_c_352_n 3.89038e-19
cc_169 N_VSS_c_163_n N_SELI_c_368_n 3.2351e-19
cc_170 N_VSS_c_175_n N_SELI_c_368_n 0.00117301f
cc_171 N_VSS_c_188_n N_SELI_c_370_n 7.32115e-19
cc_172 N_VSS_c_194_n N_SELI_c_370_n 6.85767e-19
cc_173 N_VSS_XI7.X0_PGD N_SEL_c_419_n 3.9807e-19
cc_174 N_VSS_c_171_n N_SEL_c_430_n 9.4551e-19
cc_175 N_VSS_c_194_n N_SEL_c_421_n 2.60801e-19
cc_176 N_VSS_c_188_n N_SEL_c_422_n 2.64936e-19
cc_177 N_VSS_c_155_n N_SEL_c_433_n 3.36692e-19
cc_178 N_VSS_c_171_n N_SEL_c_433_n 3.29317e-19
cc_179 N_VSS_c_185_n N_SEL_c_425_n 3.72478e-19
cc_180 N_VSS_c_155_n N_SEL_c_427_n 3.2351e-19
cc_181 N_VSS_c_171_n N_SEL_c_427_n 2.68747e-19
cc_182 N_VSS_XI7.X0_PGS N_B_XI11.X0_PGS 0.00187616f
cc_183 N_VSS_XI9.X0_PGD N_B_XI11.X0_PGS 0.00145666f
cc_184 N_VSS_c_252_p N_B_c_495_n 0.00187616f
cc_185 N_VSS_c_163_n B 3.92469e-19
cc_186 N_VSS_c_175_n B 3.5189e-19
cc_187 N_VSS_c_185_n B 2.02689e-19
cc_188 N_VSS_XI9.X0_PGD N_B_c_491_n 3.23173e-19
cc_189 N_VSS_c_147_n N_B_c_491_n 0.00295829f
cc_190 N_VSS_c_163_n N_B_c_491_n 3.5189e-19
cc_191 N_VSS_c_171_n N_B_c_491_n 6.40394e-19
cc_192 N_VSS_c_175_n N_B_c_491_n 6.81736e-19
cc_193 N_VSS_c_188_n A 2.20363e-19
cc_194 N_ZI_c_262_n N_Z_c_329_n 6.8653e-19
cc_195 N_ZI_c_271_n N_SELI_c_346_n 6.18319e-19
cc_196 N_ZI_c_277_n N_SELI_c_346_n 0.00222064f
cc_197 N_ZI_c_262_n N_SELI_c_374_n 2.5026e-19
cc_198 N_ZI_c_283_n N_SELI_c_374_n 0.00194838f
cc_199 N_ZI_c_276_n N_SELI_c_374_n 9.76295e-19
cc_200 N_ZI_c_271_n N_SELI_c_349_n 0.00164769f
cc_201 N_ZI_c_269_n N_SELI_c_350_n 0.00166258f
cc_202 N_ZI_c_277_n N_SELI_c_350_n 0.00145462f
cc_203 N_ZI_c_262_n N_SELI_c_352_n 7.59552e-19
cc_204 N_ZI_c_277_n N_SELI_c_352_n 0.00172184f
cc_205 N_ZI_c_269_n N_SELI_c_370_n 7.67117e-19
cc_206 N_ZI_c_277_n N_SELI_c_370_n 7.85627e-19
cc_207 N_ZI_c_269_n N_SELI_c_384_n 6.01706e-19
cc_208 N_ZI_c_271_n N_SELI_c_384_n 3.05282e-19
cc_209 N_ZI_c_314_p N_SELI_c_384_n 6.45182e-19
cc_210 N_ZI_c_271_n N_SELI_c_387_n 8.23018e-19
cc_211 N_ZI_c_262_n N_SEL_c_419_n 0.00374573f
cc_212 N_ZI_c_276_n N_SEL_c_439_n 4.8006e-19
cc_213 N_ZI_c_264_n N_SEL_c_420_n 9.00465e-19
cc_214 N_ZI_c_271_n N_SEL_c_420_n 0.00250758f
cc_215 N_ZI_c_277_n N_SEL_c_420_n 8.4167e-19
cc_216 N_ZI_c_269_n N_SEL_c_421_n 9.51454e-19
cc_217 N_ZI_c_271_n N_SEL_c_421_n 4.59089e-19
cc_218 N_ZI_c_314_p N_SEL_c_421_n 0.00107464f
cc_219 N_ZI_c_263_n N_SEL_c_446_n 9.00465e-19
cc_220 N_ZI_c_269_n N_SEL_c_446_n 0.00242724f
cc_221 N_ZI_c_277_n N_SEL_c_433_n 0.0014877f
cc_222 N_ZI_c_262_n N_SEL_c_427_n 5.45742e-19
cc_223 N_ZI_XI4.X0_CG N_B_XI11.X0_PGS 0.00184555f
cc_224 N_Z_c_329_n N_SELI_c_374_n 7.7787e-19
cc_225 N_Z_c_332_n N_SELI_c_374_n 0.00121421f
cc_226 N_SELI_c_343_n N_SEL_c_419_n 6.8653e-19
cc_227 N_SELI_c_346_n N_SEL_c_419_n 8.57466e-19
cc_228 N_SELI_c_349_n N_SEL_c_420_n 0.00141479f
cc_229 N_SELI_c_368_n N_SEL_c_420_n 9.76295e-19
cc_230 N_SELI_c_346_n N_SEL_c_421_n 3.66824e-19
cc_231 N_SELI_c_350_n N_SEL_c_446_n 0.00170409f
cc_232 N_SELI_c_356_n N_SEL_c_446_n 9.29204e-19
cc_233 N_SELI_c_349_n N_SEL_c_422_n 9.45347e-19
cc_234 N_SELI_c_368_n N_SEL_c_422_n 4.56568e-19
cc_235 N_SELI_c_346_n N_SEL_c_433_n 0.00216212f
cc_236 N_SELI_c_352_n N_SEL_c_433_n 7.61973e-19
cc_237 N_SELI_c_352_n N_SEL_c_425_n 0.00193122f
cc_238 N_SELI_c_350_n N_SEL_c_462_n 0.00200661f
cc_239 N_SELI_c_346_n N_SEL_c_427_n 0.00109331f
cc_240 N_SELI_c_352_n N_SEL_c_427_n 4.73568e-19
cc_241 N_SELI_c_349_n N_SEL_c_465_n 3.48267e-19
cc_242 N_SELI_c_350_n N_SEL_c_465_n 4.95293e-19
cc_243 N_SELI_c_356_n N_SEL_c_465_n 0.00480115f
cc_244 N_SELI_c_368_n N_SEL_c_465_n 9.11855e-19
cc_245 N_SELI_c_349_n N_SEL_c_428_n 4.56568e-19
cc_246 N_SELI_c_350_n N_SEL_c_428_n 3.48267e-19
cc_247 N_SELI_c_356_n N_SEL_c_428_n 9.03632e-19
cc_248 N_SELI_c_368_n N_SEL_c_428_n 0.00244546f
cc_249 N_SELI_XI11.X0_CG N_B_XI11.X0_PGS 4.83278e-19
cc_250 N_SELI_c_346_n N_B_XI11.X0_PGS 2.54355e-19
cc_251 N_SELI_c_352_n N_B_XI11.X0_PGS 8.44835e-19
cc_252 N_SELI_c_356_n N_B_XI11.X0_PGS 0.00126314f
cc_253 N_SELI_c_417_p N_A_XI10.X0_PGS 5.12461e-19
cc_254 N_SELI_c_368_n N_A_XI10.X0_PGS 0.001089f
cc_255 N_SEL_c_473_p N_B_XI11.X0_PGS 2.07014e-19
cc_256 N_SEL_c_474_p N_B_XI11.X0_PGS 4.77845e-19
cc_257 N_SEL_c_425_n N_B_XI11.X0_PGS 7.3526e-19
cc_258 N_SEL_c_427_n N_B_XI11.X0_PGS 0.00100354f
cc_259 N_SEL_c_465_n N_B_XI11.X0_PGS 0.00142122f
cc_260 N_SEL_c_462_n B 4.4727e-19
cc_261 N_SEL_c_465_n B 3.2351e-19
cc_262 N_SEL_c_462_n N_B_c_491_n 3.29317e-19
cc_263 N_SEL_c_465_n N_B_c_491_n 0.00119577f
cc_264 N_SEL_XI10.X0_CG N_A_XI10.X0_PGS 4.99479e-19
cc_265 N_SEL_c_428_n N_A_XI10.X0_PGS 0.001089f
cc_266 N_SEL_c_484_p N_A_c_537_n 9.37683e-19
cc_267 N_SEL_c_422_n A 4.54408e-19
cc_268 N_SEL_c_428_n A 3.2351e-19
cc_269 N_SEL_c_422_n N_A_c_527_n 3.2351e-19
cc_270 N_SEL_c_428_n N_A_c_527_n 2.68747e-19
cc_271 N_B_XI11.X0_PGS N_A_XI10.X0_PGS 0.00134425f
*
.ends
*
*
.subckt MUX2_HPNW8 A B S0 Y VDD VSS
xgate (VDD VSS Y S0 B A) G4_MUX2_N2
.ends
*
* File: G3_MUXI2_N2.pex.netlist
* Created: Wed Mar  9 15:09:58 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MUXI2_N2_VSS 2 4 6 8 10 12 14 29 39 51 55 60 63 68 73 78 83 92 101
+ 110 111 117 123 129 131 136 138 140 141 144 145 146 Vss
c82 146 Vss 4.28045e-19
c83 145 Vss 3.62111e-19
c84 144 Vss 3.75522e-19
c85 141 Vss 0.00260366f
c86 138 Vss 0.00496506f
c87 136 Vss 0.00156482f
c88 131 Vss 0.00130885f
c89 129 Vss 0.0025874f
c90 124 Vss 0.00128107f
c91 123 Vss 0.00657991f
c92 117 Vss 0.0039834f
c93 111 Vss 0.00549375f
c94 110 Vss 0.0044599f
c95 101 Vss 0.00833837f
c96 92 Vss 0.0039597f
c97 83 Vss 2.73987e-19
c98 78 Vss 0.00101545f
c99 73 Vss 0.00217935f
c100 68 Vss 1.35342e-19
c101 63 Vss 7.10513e-22
c102 60 Vss 0.00389683f
c103 55 Vss 0.0017936f
c104 51 Vss 0.00537538f
c105 45 Vss 0.0783825f
c106 39 Vss 0.0354115f
c107 38 Vss 0.0688416f
c108 29 Vss 0.0347733f
c109 28 Vss 0.100982f
c110 14 Vss 0.135207f
c111 10 Vss 0.135463f
c112 6 Vss 0.135561f
c113 4 Vss 0.134971f
r114 137 146 0.551426
r115 137 138 15.5878
r116 136 146 0.551426
r117 135 136 4.58464
r118 131 146 0.0828784
r119 130 145 0.494161
r120 129 138 0.652036
r121 129 130 4.41793
r122 125 145 0.128424
r123 123 135 0.652036
r124 123 124 13.0037
r125 119 124 0.652036
r126 118 144 0.494161
r127 117 145 0.494161
r128 117 118 10.2946
r129 113 144 0.128424
r130 112 140 0.326018
r131 111 144 0.494161
r132 111 112 10.1279
r133 110 140 0.326018
r134 109 141 0.14525
r135 109 110 4.54296
r136 83 131 1.82344
r137 78 101 1.16709
r138 78 125 2.16729
r139 73 119 5.2515
r140 68 92 1.16709
r141 68 113 2.16729
r142 63 141 2.334
r143 60 83 1.16709
r144 55 73 1.16709
r145 51 63 1.16709
r146 45 101 0.0476429
r147 43 45 1.8672
r148 40 43 0.0685365
r149 38 43 0.5835
r150 38 39 2.8008
r151 35 39 0.652036
r152 31 92 0.0476429
r153 29 31 1.45875
r154 28 32 0.652036
r155 28 31 1.45875
r156 25 29 0.652036
r157 14 40 3.8511
r158 12 60 0.185659
r159 10 35 3.8511
r160 8 55 0.185659
r161 6 32 3.8511
r162 4 25 3.8511
r163 2 51 0.185659
.ends

.subckt PM_G3_MUXI2_N2_VDD 2 4 6 8 10 12 14 28 38 52 56 60 62 63 66 68 72 74 75
+ 76 80 81 83 84 86 87 89 98 Vss
c93 98 Vss 0.0111581f
c94 89 Vss 0.0046197f
c95 87 Vss 4.52364e-19
c96 84 Vss 4.42749e-19
c97 83 Vss 0.0021109f
c98 81 Vss 0.00811581f
c99 80 Vss 8.64091e-19
c100 76 Vss 0.00179444f
c101 75 Vss 6.09322e-19
c102 74 Vss 0.00543501f
c103 72 Vss 0.00102525f
c104 68 Vss 0.00843754f
c105 66 Vss 0.00123499f
c106 63 Vss 6.1175e-19
c107 62 Vss 0.00356077f
c108 60 Vss 6.73464e-19
c109 56 Vss 0.00425172f
c110 52 Vss 0.00654171f
c111 44 Vss 1.28925e-19
c112 39 Vss 0.0805856f
c113 38 Vss 0.103898f
c114 29 Vss 0.0367217f
c115 28 Vss 0.101295f
c116 12 Vss 0.134871f
c117 10 Vss 0.00143442f
c118 8 Vss 0.136499f
c119 4 Vss 0.136393f
c120 2 Vss 0.13497f
r121 82 87 0.551426
r122 82 83 4.58464
r123 81 87 0.551426
r124 80 86 0.326018
r125 80 81 15.5878
r126 76 87 0.0828784
r127 76 78 1.82344
r128 74 86 0.326018
r129 74 75 10.1279
r130 72 98 1.16709
r131 70 75 0.652036
r132 70 72 2.16729
r133 69 84 0.494161
r134 68 83 0.652036
r135 68 69 13.0037
r136 64 84 0.128424
r137 64 66 5.2515
r138 62 84 0.494161
r139 62 63 7.46046
r140 60 89 1.16709
r141 58 63 0.652036
r142 58 60 2.16729
r143 56 78 1.16709
r144 52 66 1.16709
r145 44 98 0.0476429
r146 44 46 1.92555
r147 39 46 0.5835
r148 38 40 0.652036
r149 38 39 2.8008
r150 35 46 0.0685365
r151 31 89 0.0476429
r152 29 31 1.45875
r153 28 32 0.652036
r154 28 31 1.45875
r155 25 29 0.652036
r156 14 56 0.185659
r157 12 40 3.8511
r158 10 52 0.185659
r159 8 35 3.8511
r160 6 52 0.185659
r161 4 25 3.8511
r162 2 32 3.8511
.ends

.subckt PM_G3_MUXI2_N2_SELI 2 4 6 8 21 29 33 35 38 43 53 58 72 77 78 Vss
c64 78 Vss 8.06863e-19
c65 72 Vss 0.00199393f
c66 58 Vss 0.00224258f
c67 53 Vss 0.00245485f
c68 43 Vss 9.25008e-19
c69 38 Vss 0.00141078f
c70 36 Vss 0.00169592f
c71 35 Vss 0.00419199f
c72 33 Vss 0.00348196f
c73 29 Vss 0.00522942f
c74 21 Vss 0.112066f
c75 6 Vss 0.112066f
c76 4 Vss 0.00143442f
r77 77 78 0.655813
r78 76 77 3.501
r79 72 76 0.655813
r80 43 53 1.16709
r81 43 72 2.00578
r82 43 46 0.333429
r83 38 58 1.16709
r84 38 78 2.00578
r85 35 46 0.0685365
r86 35 36 7.46046
r87 31 36 0.652036
r88 31 33 7.002
r89 29 33 1.16709
r90 21 58 0.50025
r91 18 53 0.50025
r92 8 21 3.09255
r93 6 18 3.09255
r94 4 29 0.185659
r95 2 29 0.185659
.ends

.subckt PM_G3_MUXI2_N2_SEL 2 4 6 8 16 22 26 37 40 42 46 51 58 63 68 72 77 78 Vss
c64 78 Vss 7.50288e-20
c65 77 Vss 9.69437e-20
c66 72 Vss 8.26714e-19
c67 68 Vss 0.00220099f
c68 63 Vss 0.00251571f
c69 58 Vss 0.00247916f
c70 51 Vss 3.96204e-19
c71 46 Vss 8.47469e-20
c72 42 Vss 0.00123172f
c73 37 Vss 0.00197358f
c74 26 Vss 0.11221f
c75 22 Vss 0.125771f
c76 20 Vss 0.0247918f
c77 17 Vss 0.036952f
c78 16 Vss 0.188224f
c79 8 Vss 0.112066f
c80 2 Vss 0.139232f
r81 76 78 0.655813
r82 76 77 3.501
r83 72 77 0.655813
r84 54 63 1.16709
r85 54 72 2.00578
r86 51 54 0.5835
r87 49 58 1.16709
r88 46 49 0.5835
r89 42 68 1.16709
r90 42 78 2.00578
r91 38 46 0.0685365
r92 38 40 1.45875
r93 37 51 0.0685365
r94 37 40 3.12589
r95 36 58 0.0476429
r96 33 68 0.50025
r97 26 63 0.50025
r98 22 58 0.357321
r99 20 36 0.326018
r100 20 22 0.40845
r101 17 36 6.7686
r102 16 36 0.326018
r103 16 36 0.1167
r104 13 17 0.652036
r105 8 33 3.09255
r106 6 26 3.09255
r107 4 22 3.44265
r108 2 13 3.8511
.ends

.subckt PM_G3_MUXI2_N2_B 2 4 7 16 20 24 27 Vss
c24 27 Vss 0.00705011f
c25 24 Vss 6.61761e-19
c26 20 Vss 0.0287936f
c27 16 Vss 0.0658163f
c28 7 Vss 0.142266f
c29 4 Vss 0.349678f
c30 2 Vss 0.11635f
r31 24 27 1.16709
r32 16 27 0.50025
r33 16 18 1.9839
r34 12 20 0.494161
r35 9 20 0.494161
r36 8 18 0.0685365
r37 7 20 0.128424
r38 7 8 4.7847
r39 4 12 11.0281
r40 2 9 3.20925
.ends

.subckt PM_G3_MUXI2_N2_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00368622f
c33 27 Vss 0.00747653f
c34 23 Vss 0.00756091f
c35 8 Vss 0.00143442f
c36 6 Vss 0.00143442f
r37 33 35 5.91836
r38 30 33 5.08479
r39 27 35 1.16709
r40 23 30 1.16709
r41 8 27 0.185659
r42 6 23 0.185659
r43 4 27 0.185659
r44 2 23 0.185659
.ends

.subckt PM_G3_MUXI2_N2_A 2 4 14 17 23 Vss
c23 23 Vss 0.00453252f
c24 17 Vss 3.94005e-19
c25 14 Vss 0.0840432f
c26 12 Vss 1.30835e-19
c27 2 Vss 0.557463f
r28 20 23 1.16709
r29 17 20 0.0416786
r30 12 23 0.0476429
r31 12 14 1.92555
r32 7 14 0.0685365
r33 2 4 15.4044
r34 2 7 3.8511
.ends

.subckt G3_MUXI2_N2  VSS VDD SEL B Z A
*
* A	A
* Z	Z
* B	B
* SEL	SEL
* VDD	VDD
* VSS	VSS
XI6.X0 N_SELI_XI6.X0_D N_VDD_XI6.X0_PGD N_SEL_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW8
XI7.X0 N_SELI_XI7.X0_D N_VSS_XI7.X0_PGD N_SEL_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW8
XI11.X0 N_Z_XI11.X0_D N_VDD_XI11.X0_PGD N_SELI_XI11.X0_CG N_B_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW8
XI9.X0 N_Z_XI9.X0_D N_VSS_XI9.X0_PGD N_SEL_XI9.X0_CG N_B_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW8
XI10.X0 N_Z_XI10.X0_D N_VDD_XI10.X0_PGD N_SEL_XI10.X0_CG N_A_XI10.X0_PGS
+ N_VSS_XI10.X0_S TIGFET_HPNW8
XI8.X0 N_Z_XI8.X0_D N_VSS_XI8.X0_PGD N_SELI_XI8.X0_CG N_A_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW8
*
x_PM_G3_MUXI2_N2_VSS N_VSS_XI6.X0_S N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS
+ N_VSS_XI11.X0_S N_VSS_XI9.X0_PGD N_VSS_XI10.X0_S N_VSS_XI8.X0_PGD N_VSS_c_4_p
+ N_VSS_c_20_p N_VSS_c_45_p N_VSS_c_72_p N_VSS_c_27_p N_VSS_c_46_p N_VSS_c_5_p
+ N_VSS_c_26_p N_VSS_c_17_p N_VSS_c_28_p N_VSS_c_9_p N_VSS_c_19_p N_VSS_c_6_p
+ N_VSS_c_10_p N_VSS_c_11_p N_VSS_c_29_p N_VSS_c_24_p N_VSS_c_31_p N_VSS_c_34_p
+ N_VSS_c_35_p VSS N_VSS_c_50_p N_VSS_c_12_p N_VSS_c_25_p N_VSS_c_36_p Vss
+ PM_G3_MUXI2_N2_VSS
x_PM_G3_MUXI2_N2_VDD N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI7.X0_S
+ N_VDD_XI11.X0_PGD N_VDD_XI9.X0_S N_VDD_XI10.X0_PGD N_VDD_XI8.X0_S N_VDD_c_86_n
+ N_VDD_c_171_p N_VDD_c_127_p N_VDD_c_151_p N_VDD_c_87_n N_VDD_c_89_n
+ N_VDD_c_95_n N_VDD_c_96_n N_VDD_c_102_n N_VDD_c_108_n N_VDD_c_109_n
+ N_VDD_c_112_n N_VDD_c_113_n N_VDD_c_114_n N_VDD_c_115_n N_VDD_c_119_n
+ N_VDD_c_122_n VDD N_VDD_c_123_n N_VDD_c_124_n N_VDD_c_126_n Vss
+ PM_G3_MUXI2_N2_VDD
x_PM_G3_MUXI2_N2_SELI N_SELI_XI6.X0_D N_SELI_XI7.X0_D N_SELI_XI11.X0_CG
+ N_SELI_XI8.X0_CG N_SELI_c_238_p N_SELI_c_176_n N_SELI_c_178_n N_SELI_c_182_n
+ N_SELI_c_183_n N_SELI_c_197_n N_SELI_c_199_n N_SELI_c_186_n N_SELI_c_188_n
+ N_SELI_c_189_n N_SELI_c_220_p Vss PM_G3_MUXI2_N2_SELI
x_PM_G3_MUXI2_N2_SEL N_SEL_XI6.X0_CG N_SEL_XI7.X0_CG N_SEL_XI9.X0_CG
+ N_SEL_XI10.X0_CG N_SEL_c_240_n N_SEL_c_283_p N_SEL_c_284_p N_SEL_c_241_n SEL
+ N_SEL_c_242_n N_SEL_c_243_n N_SEL_c_256_n N_SEL_c_245_n N_SEL_c_271_n
+ N_SEL_c_257_n N_SEL_c_247_n N_SEL_c_249_n N_SEL_c_250_n Vss PM_G3_MUXI2_N2_SEL
x_PM_G3_MUXI2_N2_B N_B_XI11.X0_PGS N_B_XI9.X0_PGS N_B_c_304_n N_B_c_324_n
+ N_B_c_315_n B N_B_c_306_n Vss PM_G3_MUXI2_N2_B
x_PM_G3_MUXI2_N2_Z N_Z_XI11.X0_D N_Z_XI9.X0_D N_Z_XI10.X0_D N_Z_XI8.X0_D
+ N_Z_c_328_n N_Z_c_338_n N_Z_c_332_n Z Vss PM_G3_MUXI2_N2_Z
x_PM_G3_MUXI2_N2_A N_A_XI10.X0_PGS N_A_XI8.X0_PGS N_A_c_362_n A N_A_c_368_n Vss
+ PM_G3_MUXI2_N2_A
cc_1 N_VSS_XI7.X0_PGD N_VDD_XI6.X0_PGD 0.00200584f
cc_2 N_VSS_XI9.X0_PGD N_VDD_XI11.X0_PGD 2.37403e-19
cc_3 N_VSS_XI8.X0_PGD N_VDD_XI10.X0_PGD 2.37403e-19
cc_4 N_VSS_c_4_p N_VDD_c_86_n 0.00200584f
cc_5 N_VSS_c_5_p N_VDD_c_87_n 7.57561e-19
cc_6 N_VSS_c_6_p N_VDD_c_87_n 8.35657e-19
cc_7 N_VSS_c_4_p N_VDD_c_89_n 3.9313e-19
cc_8 N_VSS_c_5_p N_VDD_c_89_n 0.00161703f
cc_9 N_VSS_c_9_p N_VDD_c_89_n 2.26455e-19
cc_10 N_VSS_c_10_p N_VDD_c_89_n 0.0043279f
cc_11 N_VSS_c_11_p N_VDD_c_89_n 0.00126887f
cc_12 N_VSS_c_12_p N_VDD_c_89_n 7.74609e-19
cc_13 N_VSS_c_10_p N_VDD_c_95_n 0.00157719f
cc_14 N_VSS_XI7.X0_PGS N_VDD_c_96_n 2.59535e-19
cc_15 N_VSS_XI9.X0_PGD N_VDD_c_96_n 2.19376e-19
cc_16 N_VSS_c_5_p N_VDD_c_96_n 0.00180638f
cc_17 N_VSS_c_17_p N_VDD_c_96_n 7.4365e-19
cc_18 N_VSS_c_9_p N_VDD_c_96_n 9.55109e-19
cc_19 N_VSS_c_19_p N_VDD_c_96_n 2.70301e-19
cc_20 N_VSS_c_20_p N_VDD_c_102_n 0.00111089f
cc_21 N_VSS_c_17_p N_VDD_c_102_n 0.00161703f
cc_22 N_VSS_c_19_p N_VDD_c_102_n 2.26455e-19
cc_23 N_VSS_c_11_p N_VDD_c_102_n 0.00574413f
cc_24 N_VSS_c_24_p N_VDD_c_102_n 0.00456934f
cc_25 N_VSS_c_25_p N_VDD_c_102_n 7.61747e-19
cc_26 N_VSS_c_26_p N_VDD_c_108_n 0.00121523f
cc_27 N_VSS_c_27_p N_VDD_c_109_n 3.4118e-19
cc_28 N_VSS_c_28_p N_VDD_c_109_n 4.19648e-19
cc_29 N_VSS_c_29_p N_VDD_c_109_n 0.00755466f
cc_30 N_VSS_c_29_p N_VDD_c_112_n 0.00152669f
cc_31 N_VSS_c_31_p N_VDD_c_113_n 4.68065e-19
cc_32 N_VSS_c_29_p N_VDD_c_114_n 0.00106538f
cc_33 N_VSS_c_28_p N_VDD_c_115_n 0.00187494f
cc_34 N_VSS_c_34_p N_VDD_c_115_n 0.00339451f
cc_35 N_VSS_c_35_p N_VDD_c_115_n 0.00671233f
cc_36 N_VSS_c_36_p N_VDD_c_115_n 9.16632e-19
cc_37 N_VSS_c_17_p N_VDD_c_119_n 4.28751e-19
cc_38 N_VSS_c_19_p N_VDD_c_119_n 3.63088e-19
cc_39 N_VSS_c_35_p N_VDD_c_119_n 0.00337584f
cc_40 N_VSS_c_11_p N_VDD_c_122_n 0.0011585f
cc_41 N_VSS_c_35_p N_VDD_c_123_n 0.00100712f
cc_42 N_VSS_c_5_p N_VDD_c_124_n 3.48267e-19
cc_43 N_VSS_c_9_p N_VDD_c_124_n 6.46219e-19
cc_44 N_VSS_c_26_p N_VDD_c_126_n 2.84469e-19
cc_45 N_VSS_c_45_p N_SELI_c_176_n 3.43419e-19
cc_46 N_VSS_c_46_p N_SELI_c_176_n 3.48267e-19
cc_47 N_VSS_c_45_p N_SELI_c_178_n 3.48267e-19
cc_48 N_VSS_c_46_p N_SELI_c_178_n 5.71987e-19
cc_49 N_VSS_c_10_p N_SELI_c_178_n 2.50156e-19
cc_50 N_VSS_c_50_p N_SELI_c_178_n 2.7826e-19
cc_51 N_VSS_c_26_p N_SELI_c_182_n 0.00111908f
cc_52 N_VSS_c_17_p N_SELI_c_183_n 8.64455e-19
cc_53 N_VSS_c_19_p N_SELI_c_183_n 3.49905e-19
cc_54 N_VSS_c_35_p N_SELI_c_183_n 9.07743e-19
cc_55 N_VSS_c_17_p N_SELI_c_186_n 3.2351e-19
cc_56 N_VSS_c_19_p N_SELI_c_186_n 2.68747e-19
cc_57 N_VSS_c_29_p N_SELI_c_188_n 6.74415e-19
cc_58 N_VSS_c_35_p N_SELI_c_189_n 5.03655e-19
cc_59 N_VSS_XI7.X0_PGD N_SEL_c_240_n 4.18141e-19
cc_60 N_VSS_c_11_p N_SEL_c_241_n 5.08457e-19
cc_61 N_VSS_c_35_p N_SEL_c_242_n 7.91494e-19
cc_62 N_VSS_c_5_p N_SEL_c_243_n 5.97048e-19
cc_63 N_VSS_c_9_p N_SEL_c_243_n 3.08902e-19
cc_64 N_VSS_c_5_p N_SEL_c_245_n 3.2351e-19
cc_65 N_VSS_c_9_p N_SEL_c_245_n 2.68747e-19
cc_66 N_VSS_c_11_p N_SEL_c_247_n 0.00100236f
cc_67 N_VSS_c_29_p N_SEL_c_247_n 2.48958e-19
cc_68 N_VSS_c_35_p N_SEL_c_249_n 4.36463e-19
cc_69 N_VSS_c_29_p N_SEL_c_250_n 9.32613e-19
cc_70 N_VSS_XI7.X0_PGS N_B_c_304_n 2.56596e-19
cc_71 N_VSS_c_26_p B 0.00157463f
cc_72 N_VSS_c_72_p N_B_c_306_n 0.00246958f
cc_73 N_VSS_c_26_p N_B_c_306_n 8.835e-19
cc_74 N_VSS_c_72_p N_Z_c_328_n 3.43419e-19
cc_75 N_VSS_c_27_p N_Z_c_328_n 3.43419e-19
cc_76 N_VSS_c_26_p N_Z_c_328_n 3.48267e-19
cc_77 N_VSS_c_28_p N_Z_c_328_n 3.48267e-19
cc_78 N_VSS_c_72_p N_Z_c_332_n 3.48267e-19
cc_79 N_VSS_c_27_p N_Z_c_332_n 3.48267e-19
cc_80 N_VSS_c_26_p N_Z_c_332_n 5.71987e-19
cc_81 N_VSS_c_28_p N_Z_c_332_n 5.71987e-19
cc_82 N_VSS_c_35_p N_Z_c_332_n 6.72116e-19
cc_83 N_VDD_c_127_p N_SELI_c_176_n 3.43419e-19
cc_84 N_VDD_c_89_n N_SELI_c_176_n 3.4118e-19
cc_85 N_VDD_c_96_n N_SELI_c_176_n 3.48267e-19
cc_86 N_VDD_c_127_p N_SELI_c_178_n 3.48267e-19
cc_87 N_VDD_c_89_n N_SELI_c_178_n 4.78806e-19
cc_88 N_VDD_c_96_n N_SELI_c_178_n 7.09569e-19
cc_89 N_VDD_c_115_n N_SELI_c_183_n 6.15494e-19
cc_90 N_VDD_c_108_n N_SELI_c_197_n 4.44319e-19
cc_91 N_VDD_c_126_n N_SELI_c_197_n 3.49905e-19
cc_92 N_VDD_c_108_n N_SELI_c_199_n 3.43988e-19
cc_93 N_VDD_c_126_n N_SELI_c_199_n 2.68747e-19
cc_94 N_VDD_c_115_n N_SELI_c_186_n 3.66936e-19
cc_95 N_VDD_XI6.X0_PGD N_SEL_c_240_n 4.28909e-19
cc_96 N_VDD_c_127_p N_SEL_c_241_n 6.34806e-19
cc_97 N_VDD_c_96_n N_SEL_c_241_n 0.00105602f
cc_98 N_VDD_c_109_n N_SEL_c_242_n 2.67421e-19
cc_99 N_VDD_c_115_n N_SEL_c_242_n 6.15494e-19
cc_100 N_VDD_c_102_n N_SEL_c_256_n 2.25302e-19
cc_101 N_VDD_c_115_n N_SEL_c_257_n 3.66936e-19
cc_102 N_VDD_c_102_n N_SEL_c_247_n 4.27423e-19
cc_103 N_VDD_c_115_n N_SEL_c_249_n 2.2501e-19
cc_104 N_VDD_c_127_p N_B_c_304_n 2.2574e-19
cc_105 N_VDD_c_109_n N_Z_c_328_n 3.4118e-19
cc_106 N_VDD_c_127_p N_Z_c_338_n 3.43419e-19
cc_107 N_VDD_c_151_p N_Z_c_338_n 3.43419e-19
cc_108 N_VDD_c_96_n N_Z_c_338_n 3.48267e-19
cc_109 N_VDD_c_102_n N_Z_c_338_n 3.4118e-19
cc_110 N_VDD_c_113_n N_Z_c_338_n 3.72199e-19
cc_111 N_VDD_c_127_p N_Z_c_332_n 3.48267e-19
cc_112 N_VDD_c_151_p N_Z_c_332_n 3.48267e-19
cc_113 N_VDD_c_96_n N_Z_c_332_n 8.16241e-19
cc_114 N_VDD_c_102_n N_Z_c_332_n 4.7984e-19
cc_115 N_VDD_c_109_n N_Z_c_332_n 4.7984e-19
cc_116 N_VDD_c_113_n N_Z_c_332_n 8.08807e-19
cc_117 N_VDD_c_115_n N_Z_c_332_n 9.6188e-19
cc_118 N_VDD_XI10.X0_PGD N_A_XI10.X0_PGS 0.00151037f
cc_119 N_VDD_c_115_n N_A_XI10.X0_PGS 0.00102341f
cc_120 N_VDD_c_109_n N_A_c_362_n 3.60536e-19
cc_121 N_VDD_c_115_n N_A_c_362_n 3.92733e-19
cc_122 N_VDD_c_108_n A 5.33592e-19
cc_123 N_VDD_c_109_n A 0.00141439f
cc_124 N_VDD_c_115_n A 5.00176e-19
cc_125 N_VDD_c_126_n A 3.48267e-19
cc_126 N_VDD_XI10.X0_PGD N_A_c_368_n 3.23173e-19
cc_127 N_VDD_c_171_p N_A_c_368_n 0.00480616f
cc_128 N_VDD_c_108_n N_A_c_368_n 4.04186e-19
cc_129 N_VDD_c_109_n N_A_c_368_n 0.00120343f
cc_130 N_VDD_c_115_n N_A_c_368_n 3.66936e-19
cc_131 N_VDD_c_126_n N_A_c_368_n 6.39485e-19
cc_132 N_SELI_c_176_n N_SEL_c_240_n 6.55689e-19
cc_133 N_SELI_c_178_n N_SEL_c_240_n 9.27181e-19
cc_134 N_SELI_c_182_n N_SEL_c_240_n 4.08878e-19
cc_135 N_SELI_c_197_n N_SEL_c_241_n 0.00289751f
cc_136 N_SELI_c_183_n N_SEL_c_242_n 0.00240159f
cc_137 N_SELI_c_186_n N_SEL_c_242_n 4.99367e-19
cc_138 N_SELI_c_178_n N_SEL_c_243_n 0.0024269f
cc_139 N_SELI_c_182_n N_SEL_c_243_n 0.00289751f
cc_140 N_SELI_c_199_n N_SEL_c_256_n 5.42085e-19
cc_141 N_SELI_c_178_n N_SEL_c_245_n 0.00100994f
cc_142 N_SELI_c_182_n N_SEL_c_245_n 5.66159e-19
cc_143 N_SELI_c_199_n N_SEL_c_271_n 0.00493717f
cc_144 N_SELI_c_186_n N_SEL_c_271_n 8.7809e-19
cc_145 N_SELI_c_199_n N_SEL_c_257_n 8.69867e-19
cc_146 N_SELI_c_186_n N_SEL_c_257_n 0.00494248f
cc_147 N_SELI_c_183_n N_SEL_c_247_n 0.00165721f
cc_148 N_SELI_c_197_n N_SEL_c_247_n 4.7869e-19
cc_149 N_SELI_c_188_n N_SEL_c_247_n 9.53674e-19
cc_150 N_SELI_c_220_p N_SEL_c_247_n 7.98252e-19
cc_151 N_SELI_c_178_n N_SEL_c_249_n 3.01017e-19
cc_152 N_SELI_c_189_n N_SEL_c_249_n 0.00144491f
cc_153 N_SELI_c_197_n N_SEL_c_250_n 0.00165436f
cc_154 N_SELI_c_188_n N_SEL_c_250_n 7.97695e-19
cc_155 N_SELI_XI11.X0_CG N_B_XI11.X0_PGS 4.31731e-19
cc_156 N_SELI_c_199_n N_B_XI11.X0_PGS 6.66106e-19
cc_157 N_SELI_c_178_n N_B_XI9.X0_PGS 2.97793e-19
cc_158 N_SELI_c_182_n N_B_XI9.X0_PGS 3.99745e-19
cc_159 N_SELI_c_199_n N_B_XI9.X0_PGS 5.45575e-19
cc_160 N_SELI_c_182_n N_B_c_304_n 4.011e-19
cc_161 N_SELI_c_182_n N_B_c_315_n 5.40503e-19
cc_162 N_SELI_c_199_n N_B_c_315_n 0.00179467f
cc_163 N_SELI_c_182_n B 0.00128002f
cc_164 N_SELI_c_182_n N_B_c_306_n 0.00106912f
cc_165 N_SELI_c_178_n N_Z_c_332_n 8.31671e-19
cc_166 N_SELI_c_183_n N_Z_c_332_n 0.00208341f
cc_167 N_SELI_c_197_n N_Z_c_332_n 0.00213869f
cc_168 N_SELI_c_238_p N_A_XI10.X0_PGS 5.00154e-19
cc_169 N_SELI_c_186_n N_A_XI10.X0_PGS 0.00276355f
cc_170 N_SEL_c_283_p N_B_XI9.X0_PGS 2.04953e-19
cc_171 N_SEL_c_284_p N_B_XI9.X0_PGS 4.65537e-19
cc_172 N_SEL_c_241_n N_B_XI9.X0_PGS 8.3216e-19
cc_173 N_SEL_c_245_n N_B_XI9.X0_PGS 0.00100354f
cc_174 N_SEL_c_271_n N_B_XI9.X0_PGS 0.00202689f
cc_175 N_SEL_c_241_n N_B_c_324_n 2.88938e-19
cc_176 N_SEL_c_245_n N_B_c_324_n 7.65159e-19
cc_177 N_SEL_c_245_n N_B_c_306_n 8.68391e-19
cc_178 N_SEL_c_242_n N_Z_c_332_n 0.00189968f
cc_179 N_SEL_c_256_n N_Z_c_332_n 0.00221938f
cc_180 N_SEL_c_271_n N_Z_c_332_n 9.50991e-19
cc_181 N_SEL_c_257_n N_Z_c_332_n 9.35582e-19
cc_182 N_SEL_c_247_n N_Z_c_332_n 9.18344e-19
cc_183 N_SEL_c_249_n N_Z_c_332_n 0.0021646f
cc_184 N_SEL_c_250_n N_Z_c_332_n 9.04233e-19
cc_185 N_SEL_XI10.X0_CG N_A_XI10.X0_PGS 4.87172e-19
cc_186 N_SEL_c_257_n N_A_XI10.X0_PGS 0.00276355f
cc_187 N_SEL_c_242_n A 4.55825e-19
cc_188 N_SEL_c_257_n A 3.2351e-19
cc_189 N_SEL_c_242_n N_A_c_368_n 3.49905e-19
cc_190 N_SEL_c_257_n N_A_c_368_n 2.68747e-19
cc_191 N_B_XI11.X0_PGS N_A_XI10.X0_PGS 0.00134199f
*
.ends
*
*
.subckt MUXI2_HPNW8 A B S0 Y VDD VSS
xgate (VSS VDD S0 B Y A) G3_MUXI2_N2
.ends
*
* File: G2_NAND2_N2.pex.netlist
* Created: Fri Feb 25 16:38:49 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NAND2_N2_VSS 2 3 5 6 8 18 19 21 41 47 52 61 68 73 74 Vss
c28 74 Vss 8.01054e-19
c29 73 Vss 0.00222032f
c30 69 Vss 0.00133128f
c31 68 Vss 0.00979385f
c32 61 Vss 0.00460027f
c33 52 Vss 0.00163484f
c34 47 Vss 0.00135376f
c35 41 Vss 0.00500207f
c36 38 Vss 0.0299355f
c37 37 Vss 0.0299355f
c38 32 Vss 0.105904f
c39 26 Vss 0.0688517f
c40 21 Vss 5.38535e-20
c41 19 Vss 0.0340588f
c42 18 Vss 0.064644f
c43 8 Vss 0.138428f
c44 6 Vss 0.137392f
c45 5 Vss 0.138084f
c46 3 Vss 0.137146f
r47 73 75 0.652036
r48 73 74 4.33457
r49 66 74 0.652036
r50 66 68 7.66886
r51 65 69 0.655813
r52 65 68 8.96089
r53 52 61 1.16709
r54 52 75 2.16729
r55 47 69 1.82344
r56 41 47 1.16709
r57 33 38 0.494161
r58 32 34 0.652036
r59 32 33 2.9175
r60 28 38 0.128424
r61 27 37 0.494161
r62 26 38 0.494161
r63 26 27 2.8008
r64 22 37 0.128424
r65 21 61 0.238214
r66 19 21 1.4004
r67 18 37 0.494161
r68 18 21 1.5171
r69 15 19 0.652036
r70 8 34 3.8511
r71 6 28 3.8511
r72 5 15 3.8511
r73 3 22 3.8511
r74 2 41 0.185659
.ends

.subckt PM_G2_NAND2_N2_VDD 1 3 5 15 17 22 27 31 32 34 36 37 38 42 47 49 52 58
+ Vss
c41 58 Vss 0.00548438f
c42 50 Vss 9.22237e-19
c43 49 Vss 0.00628406f
c44 47 Vss 0.00776909f
c45 42 Vss 0.00125451f
c46 38 Vss 0.00692242f
c47 37 Vss 8.60438e-19
c48 36 Vss 0.0123084f
c49 34 Vss 0.00177187f
c50 32 Vss 8.19549e-19
c51 31 Vss 0.00243037f
c52 27 Vss 0.00484855f
c53 22 Vss 0.00385756f
c54 17 Vss 0.171989f
c55 15 Vss 0.0339269f
c56 1 Vss 0.117266f
r57 49 52 0.326018
r58 48 50 0.551426
r59 48 49 5.08479
r60 47 50 0.551426
r61 46 47 8.54411
r62 42 50 0.0828784
r63 42 44 1.82344
r64 40 58 1.16709
r65 38 46 0.655813
r66 38 40 4.37625
r67 36 52 0.326018
r68 36 37 15.6711
r69 32 34 1.76818
r70 31 37 0.652036
r71 30 32 0.657751
r72 30 31 5.04311
r73 27 44 1.16709
r74 22 34 1.16709
r75 17 58 0.428786
r76 15 17 5.3682
r77 11 15 0.652036
r78 5 27 0.185659
r79 3 22 0.185659
r80 1 11 3.1509
.ends

.subckt PM_G2_NAND2_N2_A 2 4 13 18 21 26 31 Vss
c20 31 Vss 0.00388303f
c21 26 Vss 0.00333046f
c22 18 Vss 0.00166538f
c23 13 Vss 0.112394f
c24 2 Vss 0.111896f
r25 23 31 1.16709
r26 21 23 2.54239
r27 18 26 1.16709
r28 18 21 2.83414
r29 13 31 0.50025
r30 10 26 0.50025
r31 4 13 3.09255
r32 2 10 3.09255
.ends

.subckt PM_G2_NAND2_N2_Z 2 4 6 18 22 25 28 Vss
c26 25 Vss 0.00212593f
c27 22 Vss 0.00585482f
c28 18 Vss 0.00354571f
c29 6 Vss 0.00143442f
r30 28 30 4.83471
r31 25 28 6.71025
r32 22 30 1.16709
r33 18 25 1.16709
r34 6 22 0.185659
r35 4 22 0.185659
r36 2 18 0.185659
.ends

.subckt PM_G2_NAND2_N2_B 2 4 10 11 14 18 21 Vss
c23 18 Vss 9.58314e-20
c24 14 Vss 0.181262f
c25 11 Vss 0.0357204f
c26 10 Vss 0.288966f
c27 2 Vss 0.281263f
r28 18 21 0.0416786
r29 14 18 1.16709
r30 12 14 2.1006
r31 10 12 0.652036
r32 10 11 8.92755
r33 7 11 0.652036
r34 4 14 4.3179
r35 2 7 8.57745
.ends

.subckt G2_NAND2_N2  VSS VDD A Z B
*
* B	B
* Z	Z
* A	A
* VDD	VDD
* VSS	VSS
XI12.X0 N_Z_XI12.X0_D N_VDD_XI12.X0_PGD N_A_XI12.X0_CG N_B_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW8
XI10.X0 N_Z_XI10.X0_D N_VSS_XI10.X0_PGD N_A_XI10.X0_CG N_VSS_XI10.X0_PGS
+ N_VDD_XI10.X0_S TIGFET_HPNW8
XI11.X0 N_Z_XI11.X0_D N_VSS_XI11.X0_PGD N_B_XI11.X0_CG N_VSS_XI11.X0_PGS
+ N_VDD_XI11.X0_S TIGFET_HPNW8
*
x_PM_G2_NAND2_N2_VSS N_VSS_XI12.X0_S N_VSS_XI10.X0_PGD N_VSS_XI10.X0_PGS
+ N_VSS_XI11.X0_PGD N_VSS_XI11.X0_PGS N_VSS_c_7_p N_VSS_c_8_p N_VSS_c_19_p
+ N_VSS_c_22_p N_VSS_c_6_p N_VSS_c_2_p N_VSS_c_3_p VSS N_VSS_c_11_p N_VSS_c_12_p
+ Vss PM_G2_NAND2_N2_VSS
x_PM_G2_NAND2_N2_VDD N_VDD_XI12.X0_PGD N_VDD_XI10.X0_S N_VDD_XI11.X0_S
+ N_VDD_c_62_p N_VDD_c_52_p N_VDD_c_47_p N_VDD_c_48_p N_VDD_c_29_n N_VDD_c_33_n
+ N_VDD_c_34_n N_VDD_c_35_n N_VDD_c_40_n N_VDD_c_57_p N_VDD_c_51_p N_VDD_c_59_p
+ N_VDD_c_41_n VDD N_VDD_c_45_p Vss PM_G2_NAND2_N2_VDD
x_PM_G2_NAND2_N2_A N_A_XI12.X0_CG N_A_XI10.X0_CG N_A_c_70_n N_A_c_71_n A
+ N_A_c_78_n N_A_c_74_n Vss PM_G2_NAND2_N2_A
x_PM_G2_NAND2_N2_Z N_Z_XI12.X0_D N_Z_XI10.X0_D N_Z_XI11.X0_D N_Z_c_90_n
+ N_Z_c_95_n N_Z_c_92_n Z Vss PM_G2_NAND2_N2_Z
x_PM_G2_NAND2_N2_B N_B_XI12.X0_PGS N_B_XI11.X0_CG N_B_c_116_n N_B_c_118_n
+ N_B_c_121_n N_B_c_124_n B Vss PM_G2_NAND2_N2_B
cc_1 N_VSS_XI10.X0_PGS N_VDD_c_29_n 2.7398e-19
cc_2 N_VSS_c_2_p N_VDD_c_29_n 4.50283e-19
cc_3 N_VSS_c_3_p N_VDD_c_29_n 3.70842e-19
cc_4 VSS N_VDD_c_29_n 0.00384148f
cc_5 VSS N_VDD_c_33_n 0.0016639f
cc_6 N_VSS_c_6_p N_VDD_c_34_n 4.48301e-19
cc_7 N_VSS_c_7_p N_VDD_c_35_n 0.00183557f
cc_8 N_VSS_c_8_p N_VDD_c_35_n 3.51214e-19
cc_9 N_VSS_c_2_p N_VDD_c_35_n 0.00161703f
cc_10 N_VSS_c_3_p N_VDD_c_35_n 2.03837e-19
cc_11 N_VSS_c_11_p N_VDD_c_35_n 0.00517826f
cc_12 N_VSS_c_12_p N_VDD_c_40_n 0.00104633f
cc_13 N_VSS_XI11.X0_PGS N_VDD_c_41_n 3.32059e-19
cc_14 N_VSS_c_2_p N_VDD_c_41_n 2.24202e-19
cc_15 N_VSS_c_3_p N_A_c_70_n 0.00249847f
cc_16 N_VSS_c_2_p N_A_c_71_n 2.94885e-19
cc_17 N_VSS_c_3_p N_A_c_71_n 3.71222e-19
cc_18 VSS N_A_c_71_n 0.00255481f
cc_19 N_VSS_c_19_p N_A_c_74_n 3.96531e-19
cc_20 N_VSS_c_2_p N_A_c_74_n 2.87758e-19
cc_21 N_VSS_c_3_p N_A_c_74_n 8.98435e-19
cc_22 N_VSS_c_22_p N_Z_c_90_n 3.43419e-19
cc_23 N_VSS_c_6_p N_Z_c_90_n 3.48267e-19
cc_24 N_VSS_c_6_p N_Z_c_92_n 8.92744e-19
cc_25 VSS N_Z_c_92_n 7.39325e-19
cc_26 N_VSS_XI10.X0_PGD N_B_c_116_n 8.28117e-19
cc_27 N_VSS_XI11.X0_PGD N_B_c_116_n 8.28117e-19
cc_28 N_VSS_XI10.X0_PGS N_B_c_118_n 9.94582e-19
cc_29 N_VDD_XI12.X0_PGD N_A_XI12.X0_CG 5.34714e-19
cc_30 N_VDD_XI12.X0_PGD N_A_c_78_n 2.78309e-19
cc_31 N_VDD_c_45_p N_A_c_78_n 4.44265e-19
cc_32 N_VDD_c_45_p N_Z_c_90_n 0.00132057f
cc_33 N_VDD_c_47_p N_Z_c_95_n 3.43419e-19
cc_34 N_VDD_c_48_p N_Z_c_95_n 3.43419e-19
cc_35 N_VDD_c_34_n N_Z_c_95_n 3.72199e-19
cc_36 N_VDD_c_35_n N_Z_c_95_n 3.02646e-19
cc_37 N_VDD_c_51_p N_Z_c_95_n 3.72199e-19
cc_38 N_VDD_c_52_p N_Z_c_92_n 8.40856e-19
cc_39 N_VDD_c_47_p N_Z_c_92_n 3.48267e-19
cc_40 N_VDD_c_48_p N_Z_c_92_n 3.48267e-19
cc_41 N_VDD_c_34_n N_Z_c_92_n 8.08807e-19
cc_42 N_VDD_c_35_n N_Z_c_92_n 5.981e-19
cc_43 N_VDD_c_57_p N_Z_c_92_n 0.00172841f
cc_44 N_VDD_c_51_p N_Z_c_92_n 8.49942e-19
cc_45 N_VDD_c_59_p N_Z_c_92_n 0.00179028f
cc_46 N_VDD_c_45_p N_Z_c_92_n 8.835e-19
cc_47 N_VDD_XI12.X0_PGD N_B_XI12.X0_PGS 0.00153438f
cc_48 N_VDD_c_62_p N_B_c_116_n 0.00429636f
cc_49 N_VDD_c_57_p N_B_c_121_n 2.79672e-19
cc_50 N_VDD_c_59_p N_B_c_121_n 5.52596e-19
cc_51 N_VDD_c_45_p N_B_c_121_n 7.42072e-19
cc_52 N_VDD_c_35_n N_B_c_124_n 3.13539e-19
cc_53 N_VDD_c_57_p N_B_c_124_n 3.88313e-19
cc_54 N_VDD_c_59_p N_B_c_124_n 6.60945e-19
cc_55 N_VDD_c_45_p N_B_c_124_n 2.79672e-19
cc_56 N_A_c_71_n N_Z_c_92_n 0.0082161f
cc_57 N_A_c_78_n N_Z_c_92_n 9.58524e-19
cc_58 N_A_c_74_n N_Z_c_92_n 0.00100714f
cc_59 N_A_XI12.X0_CG N_B_XI12.X0_PGS 5.00154e-19
cc_60 N_A_c_71_n N_B_XI12.X0_PGS 7.2582e-19
cc_61 N_A_c_78_n N_B_XI12.X0_PGS 5.6636e-19
cc_62 N_A_c_71_n N_B_c_116_n 3.15161e-19
cc_63 N_A_c_78_n N_B_c_116_n 7.2846e-19
cc_64 N_A_c_74_n N_B_c_116_n 0.00228839f
cc_65 N_A_c_74_n N_B_c_121_n 9.27569e-19
cc_66 N_Z_c_95_n N_B_c_116_n 3.74089e-19
cc_67 N_Z_c_92_n N_B_c_116_n 4.8079e-19
cc_68 N_Z_c_92_n N_B_c_121_n 0.00105292f
cc_69 N_Z_c_92_n N_B_c_124_n 0.00147455f
*
.ends
*
*
.subckt NAND2_HPNW8 A B Y VDD VSS
xgate (VSS VDD A Y B) G2_NAND2_N2
.ends
*
* File: G2_NOR2_N2.pex.netlist
* Created: Mon Feb 28 09:43:23 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NOR2_N2_VSS 2 4 6 18 23 28 31 36 41 50 59 60 64 65 70 77 78 80 Vss
c39 78 Vss 3.75522e-19
c40 77 Vss 0.00393043f
c41 72 Vss 0.00270228f
c42 70 Vss 0.00561311f
c43 65 Vss 8.24085e-19
c44 64 Vss 0.0017807f
c45 60 Vss 6.37548e-19
c46 59 Vss 0.00469222f
c47 50 Vss 0.0049931f
c48 41 Vss 7.10513e-22
c49 36 Vss 9.67354e-19
c50 31 Vss 0.00128167f
c51 28 Vss 0.00379689f
c52 23 Vss 0.00389355f
c53 18 Vss 0.089404f
c54 4 Vss 0.134687f
r55 77 80 0.326018
r56 76 77 4.58464
r57 72 76 0.655813
r58 71 78 0.494161
r59 70 80 0.326018
r60 70 71 10.1279
r61 66 78 0.128424
r62 64 78 0.494161
r63 64 65 4.37625
r64 59 65 0.652036
r65 58 60 0.655813
r66 58 59 15.5878
r67 41 72 1.82344
r68 36 50 1.16709
r69 36 66 2.16729
r70 31 60 1.82344
r71 28 41 1.16709
r72 23 31 1.16709
r73 16 50 0.0476429
r74 16 18 2.04225
r75 12 18 0.0685365
r76 6 28 0.185659
r77 4 12 3.8511
r78 2 23 0.185659
.ends

.subckt PM_G2_NOR2_N2_VDD 2 4 6 8 10 27 36 41 45 47 48 52 54 55 58 60 62 64 66
+ 72 78 Vss
c46 78 Vss 0.00511378f
c47 72 Vss 0.00477413f
c48 64 Vss 4.52364e-19
c49 62 Vss 0.00103884f
c50 60 Vss 6.08701e-19
c51 58 Vss 0.00137825f
c52 55 Vss 8.64106e-19
c53 54 Vss 0.00550218f
c54 52 Vss 0.00179763f
c55 49 Vss 0.00174038f
c56 48 Vss 0.00493553f
c57 47 Vss 0.00222713f
c58 45 Vss 0.00953092f
c59 41 Vss 0.00392881f
c60 37 Vss 0.129157f
c61 36 Vss 9.07184e-20
c62 27 Vss 0.035607f
c63 26 Vss 0.102409f
c64 10 Vss 0.13639f
c65 8 Vss 0.134351f
c66 4 Vss 0.13615f
c67 2 Vss 0.137207f
r68 72 75 0.05
r69 62 78 1.16709
r70 60 66 0.326018
r71 60 62 2.16729
r72 58 75 1.16709
r73 56 58 2.20896
r74 54 66 0.326018
r75 54 55 10.1696
r76 50 64 0.0828784
r77 50 52 1.82344
r78 48 56 0.652036
r79 48 49 4.37625
r80 47 55 0.652036
r81 46 64 0.551426
r82 46 47 4.58464
r83 45 64 0.551426
r84 44 49 0.652036
r85 44 45 15.5878
r86 41 52 1.16709
r87 36 72 0.0238214
r88 36 37 2.26917
r89 33 36 2.26917
r90 29 78 0.0476429
r91 27 29 1.5171
r92 26 30 0.652036
r93 26 29 1.4004
r94 23 27 0.652036
r95 20 37 0.00605528
r96 17 33 0.00605528
r97 10 30 3.8511
r98 8 23 3.8511
r99 6 41 0.185659
r100 4 17 3.8511
r101 2 20 3.8511
.ends

.subckt PM_G2_NOR2_N2_B 2 4 10 13 18 21 26 31 Vss
c20 31 Vss 0.00178268f
c21 26 Vss 0.00362926f
c22 18 Vss 0.00103738f
c23 13 Vss 0.112032f
c24 10 Vss 1.01432e-19
c25 2 Vss 0.112208f
r26 23 31 1.16709
r27 21 23 2.04225
r28 18 26 1.16709
r29 18 21 2.79246
r30 13 31 0.50025
r31 10 26 0.50025
r32 4 13 3.09255
r33 2 10 3.09255
.ends

.subckt PM_G2_NOR2_N2_Z 2 4 6 18 22 25 28 Vss
c24 25 Vss 0.00351292f
c25 22 Vss 0.00573209f
c26 18 Vss 0.00386958f
c27 6 Vss 0.00143442f
r28 28 30 4.0845
r29 25 28 6.91864
r30 22 30 1.16709
r31 18 25 1.16709
r32 6 22 0.185659
r33 4 22 0.185659
r34 2 18 0.185659
.ends

.subckt PM_G2_NOR2_N2_A 2 4 10 11 14 18 21 Vss
c17 18 Vss 2.58909e-19
c18 14 Vss 0.170846f
c19 11 Vss 0.0348505f
c20 10 Vss 0.277806f
c21 2 Vss 0.198918f
r22 18 27 1.16709
r23 18 21 0.0416786
r24 14 27 0.05
r25 12 14 1.6338
r26 10 12 0.652036
r27 10 11 8.92755
r28 7 11 0.652036
r29 4 14 4.3179
r30 2 7 5.9517
.ends

.subckt G2_NOR2_N2  VSS VDD B Z A
*
* A	A
* Z	Z
* B	B
* VDD	VDD
* VSS	VSS
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_B_XI3.X0_CG N_VDD_XI3.X0_PGS
+ N_VSS_XI3.X0_S TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VSS_XI4.X0_PGD N_B_XI4.X0_CG N_A_XI4.X0_PGS N_VDD_XI4.X0_S
+ TIGFET_HPNW8
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_VDD_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW8
*
x_PM_G2_NOR2_N2_VSS N_VSS_XI3.X0_S N_VSS_XI4.X0_PGD N_VSS_XI5.X0_S N_VSS_c_2_p
+ N_VSS_c_8_p N_VSS_c_31_p N_VSS_c_3_p N_VSS_c_6_p N_VSS_c_32_p N_VSS_c_13_p
+ N_VSS_c_4_p N_VSS_c_5_p N_VSS_c_14_p N_VSS_c_17_p N_VSS_c_15_p N_VSS_c_20_p
+ N_VSS_c_16_p VSS Vss PM_G2_NOR2_N2_VSS
x_PM_G2_NOR2_N2_VDD N_VDD_XI3.X0_PGD N_VDD_XI3.X0_PGS N_VDD_XI4.X0_S
+ N_VDD_XI5.X0_PGD N_VDD_XI5.X0_PGS N_VDD_c_41_n N_VDD_c_63_p N_VDD_c_71_p
+ N_VDD_c_42_n N_VDD_c_45_n N_VDD_c_47_n N_VDD_c_49_n N_VDD_c_50_n N_VDD_c_56_n
+ N_VDD_c_65_p N_VDD_c_57_n N_VDD_c_58_n N_VDD_c_60_n VDD N_VDD_c_66_p
+ N_VDD_c_61_n Vss PM_G2_NOR2_N2_VDD
x_PM_G2_NOR2_N2_B N_B_XI3.X0_CG N_B_XI4.X0_CG N_B_c_91_n N_B_c_102_p N_B_c_86_n
+ B N_B_c_95_n N_B_c_89_n Vss PM_G2_NOR2_N2_B
x_PM_G2_NOR2_N2_Z N_Z_XI3.X0_D N_Z_XI4.X0_D N_Z_XI5.X0_D N_Z_c_106_n N_Z_c_108_n
+ N_Z_c_110_n Z Vss PM_G2_NOR2_N2_Z
x_PM_G2_NOR2_N2_A N_A_XI4.X0_PGS N_A_XI5.X0_CG N_A_c_130_n N_A_c_133_n
+ N_A_c_135_n N_A_c_137_n A Vss PM_G2_NOR2_N2_A
cc_1 N_VSS_XI4.X0_PGD N_VDD_XI5.X0_PGD 0.00209355f
cc_2 N_VSS_c_2_p N_VDD_c_41_n 0.00209355f
cc_3 N_VSS_c_3_p N_VDD_c_42_n 0.00187494f
cc_4 N_VSS_c_4_p N_VDD_c_42_n 0.00638215f
cc_5 N_VSS_c_5_p N_VDD_c_42_n 0.00189302f
cc_6 N_VSS_c_6_p N_VDD_c_45_n 4.76491e-19
cc_7 N_VSS_c_4_p N_VDD_c_45_n 0.00344537f
cc_8 N_VSS_c_8_p N_VDD_c_47_n 3.4118e-19
cc_9 N_VSS_c_3_p N_VDD_c_47_n 9.64167e-19
cc_10 N_VSS_c_3_p N_VDD_c_49_n 4.54377e-19
cc_11 N_VSS_c_2_p N_VDD_c_50_n 3.66315e-19
cc_12 N_VSS_c_6_p N_VDD_c_50_n 0.00141228f
cc_13 N_VSS_c_13_p N_VDD_c_50_n 0.00114511f
cc_14 N_VSS_c_14_p N_VDD_c_50_n 0.00350144f
cc_15 N_VSS_c_15_p N_VDD_c_50_n 0.00445328f
cc_16 N_VSS_c_16_p N_VDD_c_50_n 7.74609e-19
cc_17 N_VSS_c_17_p N_VDD_c_56_n 0.0010632f
cc_18 N_VSS_c_15_p N_VDD_c_57_n 0.00147105f
cc_19 N_VSS_c_6_p N_VDD_c_58_n 0.00109227f
cc_20 N_VSS_c_20_p N_VDD_c_58_n 3.86251e-19
cc_21 N_VSS_c_4_p N_VDD_c_60_n 0.00116512f
cc_22 N_VSS_c_6_p N_VDD_c_61_n 3.44698e-19
cc_23 N_VSS_c_13_p N_VDD_c_61_n 6.36088e-19
cc_24 N_VSS_c_6_p N_B_c_86_n 5.58916e-19
cc_25 N_VSS_c_13_p N_B_c_86_n 3.52408e-19
cc_26 N_VSS_c_4_p N_B_c_86_n 0.00152314f
cc_27 N_VSS_c_6_p N_B_c_89_n 3.2351e-19
cc_28 N_VSS_c_13_p N_B_c_89_n 0.00119577f
cc_29 N_VSS_c_8_p N_Z_c_106_n 3.43419e-19
cc_30 N_VSS_c_3_p N_Z_c_106_n 3.48267e-19
cc_31 N_VSS_c_31_p N_Z_c_108_n 3.43419e-19
cc_32 N_VSS_c_32_p N_Z_c_108_n 3.48267e-19
cc_33 N_VSS_c_8_p N_Z_c_110_n 3.48267e-19
cc_34 N_VSS_c_31_p N_Z_c_110_n 3.48267e-19
cc_35 N_VSS_c_3_p N_Z_c_110_n 8.54909e-19
cc_36 N_VSS_c_32_p N_Z_c_110_n 5.71987e-19
cc_37 N_VSS_c_4_p N_Z_c_110_n 7.7813e-19
cc_38 N_VSS_c_15_p N_Z_c_110_n 2.40801e-19
cc_39 N_VSS_XI4.X0_PGD N_A_c_130_n 9.55607e-19
cc_40 N_VDD_c_63_p N_B_c_91_n 8.8401e-19
cc_41 N_VDD_c_42_n N_B_c_86_n 0.00264899f
cc_42 N_VDD_c_65_p N_B_c_86_n 5.00177e-19
cc_43 N_VDD_c_66_p N_B_c_86_n 3.55951e-19
cc_44 N_VDD_c_42_n N_B_c_95_n 5.06499e-19
cc_45 N_VDD_c_65_p N_B_c_95_n 3.43988e-19
cc_46 N_VDD_c_66_p N_B_c_95_n 2.75266e-19
cc_47 N_VDD_c_42_n N_B_c_89_n 3.66936e-19
cc_48 N_VDD_c_71_p N_Z_c_108_n 3.43419e-19
cc_49 N_VDD_c_49_n N_Z_c_108_n 3.72199e-19
cc_50 N_VDD_c_50_n N_Z_c_108_n 3.4118e-19
cc_51 N_VDD_c_71_p N_Z_c_110_n 3.48267e-19
cc_52 N_VDD_c_42_n N_Z_c_110_n 9.15147e-19
cc_53 N_VDD_c_49_n N_Z_c_110_n 7.92786e-19
cc_54 N_VDD_c_50_n N_Z_c_110_n 4.80596e-19
cc_55 N_VDD_XI3.X0_PGD N_A_c_130_n 5.1398e-19
cc_56 N_VDD_XI5.X0_PGD N_A_c_130_n 2.51476e-19
cc_57 N_VDD_XI3.X0_PGS N_A_c_133_n 6.75208e-19
cc_58 N_VDD_c_42_n N_A_c_133_n 4.39208e-19
cc_59 N_VDD_c_58_n N_A_c_135_n 3.47446e-19
cc_60 N_VDD_c_61_n N_A_c_135_n 0.00119807f
cc_61 N_VDD_c_58_n N_A_c_137_n 4.24105e-19
cc_62 N_VDD_c_61_n N_A_c_137_n 3.26762e-19
cc_63 N_B_c_86_n N_Z_c_110_n 0.00741085f
cc_64 N_B_c_95_n N_Z_c_110_n 0.0010409f
cc_65 N_B_c_89_n N_Z_c_110_n 9.42705e-19
cc_66 N_B_c_102_p N_A_XI4.X0_PGS 5.00154e-19
cc_67 N_B_c_89_n N_A_XI4.X0_PGS 7.86826e-19
cc_68 N_B_c_95_n N_A_c_130_n 0.00159105f
cc_69 N_B_c_89_n N_A_c_135_n 7.50183e-19
cc_70 N_Z_c_108_n N_A_c_130_n 4.45882e-19
cc_71 N_Z_c_110_n N_A_c_130_n 9.61158e-19
cc_72 N_Z_c_110_n N_A_c_135_n 0.00108982f
cc_73 N_Z_c_110_n N_A_c_137_n 0.00155484f
*
.ends
*
*
.subckt NOR2_HPNW8 A B Y VDD VSS
xgate (VSS VDD B Y A) G2_NOR2_N2
.ends
*
* File: G2_OAI21_N2.pex.netlist
* Created: Wed Mar  2 11:29:59 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_OAI21_N2_VSS 2 4 6 8 10 22 29 37 42 45 50 55 64 73 74 78 84 86 91
+ 94 Vss
c51 92 Vss 5.73928e-19
c52 91 Vss 0.00804514f
c53 86 Vss 0.00176984f
c54 84 Vss 0.00284334f
c55 79 Vss 0.00136792f
c56 78 Vss 0.00717474f
c57 74 Vss 6.26507e-19
c58 73 Vss 0.00636709f
c59 64 Vss 0.0055272f
c60 55 Vss 2.73987e-19
c61 50 Vss 0.00176484f
c62 45 Vss 0.00142483f
c63 42 Vss 0.00389683f
c64 37 Vss 0.00480057f
c65 33 Vss 0.0307649f
c66 29 Vss 6.10339e-20
c67 26 Vss 0.101243f
c68 22 Vss 0.0345703f
c69 21 Vss 0.0712517f
c70 10 Vss 0.136616f
c71 8 Vss 0.135636f
c72 4 Vss 0.135245f
r73 91 94 0.326018
r74 90 91 16.0879
r75 86 90 0.655813
r76 85 92 0.494161
r77 84 94 0.326018
r78 84 85 4.33457
r79 80 92 0.128424
r80 78 92 0.494161
r81 78 79 10.1696
r82 73 79 0.652036
r83 72 74 0.655813
r84 72 73 16.0879
r85 55 86 1.82344
r86 50 64 1.16709
r87 50 80 2.16729
r88 45 74 1.82344
r89 42 55 1.16709
r90 37 45 1.16709
r91 29 64 0.238214
r92 27 33 0.494161
r93 27 29 1.5171
r94 26 30 0.652036
r95 26 29 1.4004
r96 23 33 0.128424
r97 21 33 0.494161
r98 21 22 2.8008
r99 18 22 0.652036
r100 10 30 3.8511
r101 8 23 3.8511
r102 6 42 0.185659
r103 4 18 3.8511
r104 2 37 0.185659
.ends

.subckt PM_G2_OAI21_N2_VDD 2 4 6 8 30 35 38 39 41 43 47 49 51 56 59 65 Vss
c49 65 Vss 0.00587512f
c50 57 Vss 5.34798e-19
c51 56 Vss 0.0102152f
c52 55 Vss 0.00177964f
c53 51 Vss 0.00246273f
c54 49 Vss 0.00378116f
c55 47 Vss 0.00135688f
c56 43 Vss 0.00167028f
c57 41 Vss 8.22855e-19
c58 40 Vss 0.00177964f
c59 39 Vss 0.00981195f
c60 38 Vss 0.0104045f
c61 35 Vss 0.0039168f
c62 30 Vss 0.00399277f
c63 25 Vss 0.0856551f
c64 19 Vss 0.0340946f
c65 18 Vss 0.0688517f
c66 6 Vss 0.137594f
c67 2 Vss 0.137999f
r68 55 59 0.326018
r69 55 56 16.0879
r70 51 56 0.655813
r71 51 53 1.82344
r72 50 57 0.494161
r73 49 59 0.326018
r74 49 50 4.37625
r75 47 65 1.16709
r76 45 57 0.128424
r77 45 47 2.16729
r78 41 43 1.82344
r79 39 57 0.494161
r80 39 40 10.1279
r81 38 41 0.655813
r82 37 40 0.652036
r83 37 38 16.0879
r84 35 53 1.16709
r85 30 43 1.16709
r86 25 65 0.238214
r87 23 25 2.04225
r88 20 23 0.0685365
r89 18 23 0.5835
r90 18 19 2.8008
r91 15 19 0.652036
r92 8 35 0.185659
r93 6 20 3.8511
r94 4 30 0.185659
r95 2 15 3.8511
.ends

.subckt PM_G2_OAI21_N2_B 2 4 13 18 21 26 31 Vss
c21 31 Vss 0.00395418f
c22 26 Vss 0.00337806f
c23 18 Vss 6.82306e-19
c24 13 Vss 0.113634f
c25 10 Vss 1.97908e-19
c26 2 Vss 0.112205f
r27 23 31 1.16709
r28 21 23 1.7505
r29 18 26 1.16709
r30 18 21 3.08421
r31 13 31 0.476429
r32 10 26 0.50025
r33 4 13 3.1509
r34 2 10 3.09255
.ends

.subckt PM_G2_OAI21_N2_A 2 4 13 18 21 26 31 36 44 46 Vss
c41 46 Vss 1.69877e-19
c42 36 Vss 0.00272497f
c43 31 Vss 0.00729791f
c44 26 Vss 0.0034552f
c45 21 Vss 0.00215165f
c46 18 Vss 0.0860045f
c47 13 Vss 5.54498e-20
c48 4 Vss 0.112066f
c49 2 Vss 0.138617f
r50 40 46 0.655813
r51 26 36 1.16709
r52 26 46 4.52212
r53 21 31 1.16709
r54 21 44 0.0416786
r55 21 40 10.8364
r56 18 31 0.238214
r57 15 18 1.92555
r58 13 36 0.50025
r59 7 15 0.0685365
r60 4 13 3.09255
r61 2 7 3.8511
.ends

.subckt PM_G2_OAI21_N2_Z 2 4 6 8 23 27 30 33 Vss
c33 30 Vss 0.0014926f
c34 27 Vss 0.00690919f
c35 23 Vss 0.00596354f
c36 8 Vss 0.00143442f
c37 6 Vss 0.00143442f
r38 33 35 4.20954
r39 30 33 6.79361
r40 27 35 1.16709
r41 23 30 1.16709
r42 8 27 0.185659
r43 6 23 0.185659
r44 4 27 0.185659
r45 2 23 0.185659
.ends

.subckt PM_G2_OAI21_N2_C 2 4 6 13 14 17 24 27 30 Vss
c31 27 Vss 4.25339e-19
c32 24 Vss 0.0812712f
c33 17 Vss 0.202681f
c34 14 Vss 0.0348616f
c35 13 Vss 0.246708f
c36 4 Vss 0.235568f
c37 2 Vss 0.235767f
r38 27 30 0.0833571
r39 23 24 2.04225
r40 20 24 0.0685365
r41 17 27 1.16709
r42 15 23 0.0685365
r43 15 17 2.8008
r44 13 23 0.5835
r45 13 14 8.92755
r46 10 14 0.652036
r47 6 17 4.3179
r48 4 20 7.1187
r49 2 10 7.1187
.ends

.subckt G2_OAI21_N2  VSS VDD B A Z C
*
* C	C
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_B_XI3.X0_CG N_C_XI3.X0_PGS N_VSS_XI3.X0_S
+ TIGFET_HPNW8
XI0.X0 N_Z_XI0.X0_D N_VSS_XI0.X0_PGD N_B_XI0.X0_CG N_A_XI0.X0_PGS N_VDD_XI0.X0_S
+ TIGFET_HPNW8
XI4.X0 N_Z_XI4.X0_D N_VDD_XI4.X0_PGD N_A_XI4.X0_CG N_C_XI4.X0_PGS N_VSS_XI4.X0_S
+ TIGFET_HPNW8
XI2.X0 N_Z_XI2.X0_D N_VSS_XI2.X0_PGD N_C_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW8
*
x_PM_G2_OAI21_N2_VSS N_VSS_XI3.X0_S N_VSS_XI0.X0_PGD N_VSS_XI4.X0_S
+ N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS N_VSS_c_29_p N_VSS_c_46_p N_VSS_c_1_p
+ N_VSS_c_9_p N_VSS_c_2_p N_VSS_c_21_p N_VSS_c_10_p N_VSS_c_22_p N_VSS_c_3_p
+ N_VSS_c_4_p N_VSS_c_8_p N_VSS_c_12_p N_VSS_c_11_p N_VSS_c_14_p VSS Vss
+ PM_G2_OAI21_N2_VSS
x_PM_G2_OAI21_N2_VDD N_VDD_XI3.X0_PGD N_VDD_XI0.X0_S N_VDD_XI4.X0_PGD
+ N_VDD_XI2.X0_S N_VDD_c_84_p N_VDD_c_85_p N_VDD_c_52_n N_VDD_c_56_n
+ N_VDD_c_57_n N_VDD_c_58_n N_VDD_c_77_p N_VDD_c_60_n N_VDD_c_63_n N_VDD_c_66_n
+ VDD N_VDD_c_74_p Vss PM_G2_OAI21_N2_VDD
x_PM_G2_OAI21_N2_B N_B_XI3.X0_CG N_B_XI0.X0_CG N_B_c_109_p N_B_c_101_n B
+ N_B_c_104_n N_B_c_105_n Vss PM_G2_OAI21_N2_B
x_PM_G2_OAI21_N2_A N_A_XI0.X0_PGS N_A_XI4.X0_CG N_A_c_137_n N_A_c_145_n
+ N_A_c_123_n N_A_c_128_n N_A_c_130_n N_A_c_134_n A N_A_c_135_n Vss
+ PM_G2_OAI21_N2_A
x_PM_G2_OAI21_N2_Z N_Z_XI3.X0_D N_Z_XI0.X0_D N_Z_XI4.X0_D N_Z_XI2.X0_D
+ N_Z_c_163_n N_Z_c_174_n N_Z_c_167_n Z Vss PM_G2_OAI21_N2_Z
x_PM_G2_OAI21_N2_C N_C_XI3.X0_PGS N_C_XI4.X0_PGS N_C_XI2.X0_CG N_C_c_196_n
+ N_C_c_218_n N_C_c_198_n N_C_c_201_n N_C_c_202_n C Vss PM_G2_OAI21_N2_C
cc_1 N_VSS_c_1_p N_VDD_c_52_n 9.5668e-19
cc_2 N_VSS_c_2_p N_VDD_c_52_n 0.00165395f
cc_3 N_VSS_c_3_p N_VDD_c_52_n 0.00691557f
cc_4 N_VSS_c_4_p N_VDD_c_52_n 0.00189413f
cc_5 N_VSS_c_2_p N_VDD_c_56_n 9.07068e-19
cc_6 N_VSS_c_3_p N_VDD_c_57_n 0.0016897f
cc_7 N_VSS_c_2_p N_VDD_c_58_n 4.55601e-19
cc_8 N_VSS_c_8_p N_VDD_c_58_n 4.44911e-19
cc_9 N_VSS_c_9_p N_VDD_c_60_n 3.02646e-19
cc_10 N_VSS_c_10_p N_VDD_c_60_n 4.09912e-19
cc_11 N_VSS_c_11_p N_VDD_c_60_n 4.66923e-19
cc_12 N_VSS_c_12_p N_VDD_c_63_n 4.44911e-19
cc_13 N_VSS_c_11_p N_VDD_c_63_n 4.55601e-19
cc_14 N_VSS_c_14_p N_VDD_c_63_n 0.00176782f
cc_15 N_VSS_c_9_p N_VDD_c_66_n 9.5668e-19
cc_16 N_VSS_c_10_p N_VDD_c_66_n 0.00165395f
cc_17 N_VSS_c_11_p N_VDD_c_66_n 0.00189413f
cc_18 N_VSS_c_14_p N_VDD_c_66_n 0.00744813f
cc_19 N_VSS_c_3_p N_B_c_101_n 5.69535e-19
cc_20 N_VSS_XI0.X0_PGD N_A_XI0.X0_PGS 0.00176902f
cc_21 N_VSS_c_21_p N_A_c_123_n 8.59446e-19
cc_22 N_VSS_c_22_p N_A_c_123_n 3.44698e-19
cc_23 N_VSS_c_3_p N_A_c_123_n 0.003788f
cc_24 N_VSS_c_8_p N_A_c_123_n 0.00211252f
cc_25 N_VSS_c_14_p N_A_c_123_n 0.00180094f
cc_26 N_VSS_c_8_p N_A_c_128_n 7.40806e-19
cc_27 N_VSS_c_14_p N_A_c_128_n 7.9739e-19
cc_28 N_VSS_XI0.X0_PGD N_A_c_130_n 3.11814e-19
cc_29 N_VSS_c_29_p N_A_c_130_n 0.00322564f
cc_30 N_VSS_c_21_p N_A_c_130_n 3.44698e-19
cc_31 N_VSS_c_22_p N_A_c_130_n 6.61253e-19
cc_32 N_VSS_c_22_p N_A_c_134_n 2.86526e-19
cc_33 N_VSS_c_3_p N_A_c_135_n 0.00310102f
cc_34 N_VSS_c_1_p N_Z_c_163_n 3.43419e-19
cc_35 N_VSS_c_9_p N_Z_c_163_n 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_c_163_n 3.48267e-19
cc_37 N_VSS_c_10_p N_Z_c_163_n 3.48267e-19
cc_38 N_VSS_c_1_p N_Z_c_167_n 3.48267e-19
cc_39 N_VSS_c_9_p N_Z_c_167_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_167_n 5.71987e-19
cc_41 N_VSS_c_10_p N_Z_c_167_n 5.71987e-19
cc_42 N_VSS_c_8_p N_Z_c_167_n 3.27942e-19
cc_43 N_VSS_c_14_p N_Z_c_167_n 6.37542e-19
cc_44 N_VSS_XI0.X0_PGD N_C_c_196_n 6.82193e-19
cc_45 N_VSS_XI2.X0_PGD N_C_c_196_n 6.82193e-19
cc_46 N_VSS_c_46_p N_C_c_198_n 4.58946e-19
cc_47 N_VSS_c_21_p N_C_c_198_n 2.87758e-19
cc_48 N_VSS_c_22_p N_C_c_198_n 0.00236077f
cc_49 N_VSS_XI2.X0_PGS N_C_c_201_n 8.15793e-19
cc_50 N_VSS_c_21_p N_C_c_202_n 2.83343e-19
cc_51 N_VSS_c_22_p N_C_c_202_n 2.87758e-19
cc_52 N_VDD_c_52_n N_B_c_101_n 0.00231792f
cc_53 N_VDD_c_56_n N_B_c_101_n 2.08521e-19
cc_54 N_VDD_c_52_n N_B_c_104_n 3.66936e-19
cc_55 N_VDD_c_52_n N_B_c_105_n 4.5927e-19
cc_56 N_VDD_c_74_p N_A_XI4.X0_CG 0.00253477f
cc_57 N_VDD_c_74_p N_A_c_137_n 6.39343e-19
cc_58 N_VDD_c_56_n N_A_c_128_n 7.76297e-19
cc_59 N_VDD_c_77_p N_A_c_128_n 5.10019e-19
cc_60 N_VDD_c_66_n N_A_c_128_n 6.23587e-19
cc_61 N_VDD_c_74_p N_A_c_128_n 3.18657e-19
cc_62 N_VDD_c_66_n N_A_c_134_n 3.66936e-19
cc_63 N_VDD_c_74_p N_A_c_134_n 6.82215e-19
cc_64 N_VDD_c_52_n N_A_c_135_n 6.11072e-19
cc_65 N_VDD_c_56_n N_Z_c_163_n 3.02646e-19
cc_66 N_VDD_c_84_p N_Z_c_174_n 3.43419e-19
cc_67 N_VDD_c_85_p N_Z_c_174_n 3.43419e-19
cc_68 N_VDD_c_58_n N_Z_c_174_n 3.72199e-19
cc_69 N_VDD_c_63_n N_Z_c_174_n 3.72199e-19
cc_70 N_VDD_c_84_p N_Z_c_167_n 3.48267e-19
cc_71 N_VDD_c_85_p N_Z_c_167_n 3.48267e-19
cc_72 N_VDD_c_52_n N_Z_c_167_n 7.99049e-19
cc_73 N_VDD_c_56_n N_Z_c_167_n 6.12187e-19
cc_74 N_VDD_c_58_n N_Z_c_167_n 5.09542e-19
cc_75 N_VDD_c_63_n N_Z_c_167_n 7.72285e-19
cc_76 N_VDD_c_66_n N_Z_c_167_n 0.00141871f
cc_77 N_VDD_c_52_n N_C_XI3.X0_PGS 6.13097e-19
cc_78 N_VDD_c_66_n N_C_XI4.X0_PGS 6.32546e-19
cc_79 N_VDD_XI3.X0_PGD N_C_c_196_n 6.82193e-19
cc_80 N_VDD_XI4.X0_PGD N_C_c_196_n 6.82193e-19
cc_81 N_VDD_c_66_n N_C_c_198_n 5.55044e-19
cc_82 N_VDD_c_66_n N_C_c_202_n 5.04211e-19
cc_83 N_B_c_105_n N_A_c_145_n 4.64013e-19
cc_84 N_B_c_101_n N_A_c_123_n 0.0028587f
cc_85 N_B_c_105_n N_A_c_123_n 2.87758e-19
cc_86 N_B_c_109_p N_A_c_130_n 0.00249847f
cc_87 N_B_c_101_n N_A_c_130_n 3.4348e-19
cc_88 N_B_c_105_n N_A_c_130_n 6.82215e-19
cc_89 N_B_c_104_n N_A_c_134_n 8.86454e-19
cc_90 N_B_c_101_n N_A_c_135_n 7.33011e-19
cc_91 N_B_c_101_n N_Z_c_167_n 0.00671f
cc_92 N_B_c_104_n N_Z_c_167_n 9.58174e-19
cc_93 N_B_c_105_n N_Z_c_167_n 0.00100281f
cc_94 N_B_XI3.X0_CG N_C_XI3.X0_PGS 4.87172e-19
cc_95 N_B_c_104_n N_C_XI3.X0_PGS 0.001089f
cc_96 N_B_c_104_n N_C_c_196_n 6.02551e-19
cc_97 N_B_c_105_n N_C_c_196_n 0.00129343f
cc_98 N_B_c_105_n N_C_c_198_n 9.54365e-19
cc_99 N_A_c_123_n N_Z_c_167_n 0.00174866f
cc_100 N_A_c_128_n N_Z_c_167_n 0.00351012f
cc_101 N_A_c_134_n N_Z_c_167_n 9.53427e-19
cc_102 N_A_XI4.X0_CG N_C_XI4.X0_PGS 4.87172e-19
cc_103 N_A_c_134_n N_C_XI4.X0_PGS 0.001089f
cc_104 N_A_c_134_n N_C_c_196_n 0.00151445f
cc_105 N_A_XI0.X0_PGS N_C_c_218_n 8.15793e-19
cc_106 N_A_c_128_n N_C_c_198_n 5.38228e-19
cc_107 N_A_c_134_n N_C_c_198_n 0.00209031f
cc_108 N_A_c_128_n N_C_c_202_n 8.16123e-19
cc_109 N_Z_c_163_n N_C_c_196_n 3.50149e-19
cc_110 N_Z_c_174_n N_C_c_196_n 3.50149e-19
cc_111 N_Z_c_167_n N_C_c_196_n 3.56555e-19
cc_112 N_Z_c_167_n N_C_c_198_n 0.00102535f
cc_113 N_Z_c_167_n N_C_c_202_n 0.00141616f
*
.ends
*
*
.subckt OAI21_HPNW8 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 A0 Y B0) G2_OAI21_N2
.ends
*
* File: G3_OR2_N2.pex.netlist
* Created: Tue Mar  1 12:00:05 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_OR2_N2_VSS 2 4 6 8 10 12 28 29 38 44 49 52 57 62 67 76 85 90 91 93
+ 97 98 103 109 115 116 Vss
c69 116 Vss 3.88979e-19
c70 115 Vss 3.75522e-19
c71 109 Vss 0.00356171f
c72 103 Vss 0.00288176f
c73 98 Vss 8.31407e-19
c74 97 Vss 0.0017807f
c75 91 Vss 6.38539e-19
c76 90 Vss 0.00489715f
c77 85 Vss 0.00399322f
c78 76 Vss 0.00493786f
c79 67 Vss 5.89061e-19
c80 62 Vss 7.90818e-19
c81 57 Vss 8.66334e-19
c82 52 Vss 0.00128155f
c83 49 Vss 0.00709351f
c84 44 Vss 0.00389355f
c85 38 Vss 0.0895618f
c86 29 Vss 0.0349332f
c87 28 Vss 0.0997249f
c88 12 Vss 0.134814f
c89 10 Vss 0.13405f
c90 8 Vss 0.00143442f
c91 4 Vss 0.134687f
r92 110 116 0.494161
r93 109 111 0.652036
r94 109 110 7.46046
r95 105 116 0.128424
r96 104 115 0.494161
r97 103 116 0.494161
r98 103 104 7.46046
r99 99 115 0.128424
r100 97 115 0.494161
r101 97 98 4.37625
r102 91 93 0.765844
r103 90 98 0.652036
r104 89 91 0.655813
r105 89 90 15.5878
r106 67 85 1.16709
r107 67 111 2.16729
r108 62 105 5.2515
r109 57 76 1.16709
r110 57 99 2.16729
r111 52 93 1.05759
r112 49 62 1.16709
r113 44 52 1.16709
r114 36 76 0.0476429
r115 36 38 2.04225
r116 31 85 0.0476429
r117 29 31 1.45875
r118 28 32 0.652036
r119 28 31 1.45875
r120 25 29 0.652036
r121 22 38 0.0685365
r122 12 32 3.8511
r123 10 25 3.8511
r124 8 49 0.185659
r125 6 49 0.185659
r126 4 22 3.8511
r127 2 44 0.185659
.ends

.subckt PM_G3_OR2_N2_VDD 2 4 6 8 10 12 14 16 37 46 56 62 67 70 72 73 77 79 80 83
+ 87 89 93 95 97 102 104 105 106 107 113 119 124 Vss
c78 124 Vss 0.00436477f
c79 119 Vss 0.00478009f
c80 113 Vss 0.00477414f
c81 107 Vss 2.39889e-19
c82 106 Vss 2.39889e-19
c83 105 Vss 4.52364e-19
c84 102 Vss 0.00334204f
c85 97 Vss 0.00329381f
c86 95 Vss 0.00842218f
c87 93 Vss 5.48147e-19
c88 89 Vss 0.00206676f
c89 87 Vss 4.88586e-19
c90 83 Vss 0.00135406f
c91 80 Vss 8.68155e-19
c92 79 Vss 0.00563376f
c93 77 Vss 0.0017975f
c94 73 Vss 0.0049339f
c95 72 Vss 0.00221679f
c96 70 Vss 0.00947695f
c97 69 Vss 0.00174028f
c98 67 Vss 0.00532741f
c99 62 Vss 0.00393183f
c100 57 Vss 0.129157f
c101 56 Vss 9.10906e-20
c102 47 Vss 0.0358563f
c103 46 Vss 0.101295f
c104 37 Vss 0.035607f
c105 36 Vss 0.101546f
c106 14 Vss 0.134527f
c107 12 Vss 0.134502f
c108 10 Vss 0.13477f
c109 8 Vss 0.134351f
c110 4 Vss 0.136655f
c111 2 Vss 0.137748f
r112 113 116 0.05
r113 101 102 4.58464
r114 97 101 0.655813
r115 97 99 1.82344
r116 96 107 0.494161
r117 95 102 0.652036
r118 95 96 10.1279
r119 93 124 1.16709
r120 91 107 0.128424
r121 91 93 2.16729
r122 90 106 0.494161
r123 89 107 0.494161
r124 89 90 4.54296
r125 87 119 1.16709
r126 85 106 0.128424
r127 85 87 2.16729
r128 83 116 1.16709
r129 81 83 2.16729
r130 79 106 0.494161
r131 79 80 10.1696
r132 75 105 0.0828784
r133 75 77 1.82344
r134 74 104 0.326018
r135 73 81 0.652036
r136 73 74 4.37625
r137 72 80 0.652036
r138 71 105 0.551426
r139 71 72 4.58464
r140 70 105 0.551426
r141 69 104 0.326018
r142 69 70 15.5461
r143 67 99 1.16709
r144 62 77 1.16709
r145 56 113 0.0238214
r146 56 57 2.26917
r147 53 56 2.26917
r148 49 124 0.0476429
r149 47 49 1.45875
r150 46 50 0.652036
r151 46 49 1.45875
r152 43 47 0.652036
r153 39 119 0.0476429
r154 37 39 1.5171
r155 36 40 0.652036
r156 36 39 1.4004
r157 33 37 0.652036
r158 30 57 0.00605528
r159 27 53 0.00605528
r160 16 67 0.185659
r161 14 43 3.8511
r162 12 50 3.8511
r163 10 40 3.8511
r164 8 33 3.8511
r165 6 62 0.185659
r166 4 27 3.8511
r167 2 30 3.8511
.ends

.subckt PM_G3_OR2_N2_B 2 4 10 13 18 21 26 31 Vss
c21 31 Vss 0.00178268f
c22 26 Vss 0.00362926f
c23 18 Vss 9.47382e-19
c24 13 Vss 0.112032f
c25 10 Vss 1.01848e-19
c26 2 Vss 0.112208f
r27 23 31 1.16709
r28 21 23 2.20896
r29 18 26 1.16709
r30 18 21 2.62575
r31 13 31 0.50025
r32 10 26 0.50025
r33 4 13 3.09255
r34 2 10 3.09255
.ends

.subckt PM_G3_OR2_N2_NET21 2 4 6 8 10 24 27 38 42 45 53 66 70 Vss
c39 70 Vss 0.00743392f
c40 66 Vss 0.0057739f
c41 53 Vss 0.00155523f
c42 45 Vss 0.00308587f
c43 42 Vss 0.00569159f
c44 38 Vss 0.00386958f
c45 27 Vss 1.05421e-19
c46 24 Vss 0.225855f
c47 21 Vss 0.125908f
c48 19 Vss 0.0247918f
c49 10 Vss 0.139046f
c50 6 Vss 0.00143442f
r51 70 74 0.655813
r52 53 66 1.16709
r53 53 74 2.08393
r54 48 70 7.03847
r55 48 50 5.835
r56 45 48 5.16814
r57 42 50 1.16709
r58 38 45 1.16709
r59 27 66 0.0476429
r60 25 27 0.326018
r61 25 27 0.1167
r62 24 28 0.652036
r63 24 27 6.7686
r64 21 66 0.357321
r65 19 27 0.326018
r66 19 21 0.40845
r67 10 28 3.8511
r68 8 21 3.44265
r69 6 42 0.185659
r70 4 42 0.185659
r71 2 38 0.185659
.ends

.subckt PM_G3_OR2_N2_A 2 4 10 11 14 18 21 Vss
c21 18 Vss 3.18373e-19
c22 14 Vss 0.170625f
c23 11 Vss 0.0348505f
c24 10 Vss 0.277805f
c25 2 Vss 0.198918f
r26 18 27 1.16709
r27 18 21 0.0833571
r28 14 27 0.05
r29 12 14 1.6338
r30 10 12 0.652036
r31 10 11 8.92755
r32 7 11 0.652036
r33 4 14 4.3179
r34 2 7 5.9517
.ends

.subckt PM_G3_OR2_N2_Z 2 4 13 16 19 Vss
c12 13 Vss 0.00522942f
c13 4 Vss 0.00143442f
r14 16 19 0.0353636
r15 13 19 1.16709
r16 4 13 0.185659
r17 2 13 0.185659
.ends

.subckt G3_OR2_N2  VSS VDD B A Z
*
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI7.X0 N_NET21_XI7.X0_D N_VDD_XI7.X0_PGD N_B_XI7.X0_CG N_VDD_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW8
XI5.X0 N_NET21_XI5.X0_D N_VSS_XI5.X0_PGD N_B_XI5.X0_CG N_A_XI5.X0_PGS
+ N_VDD_XI5.X0_S TIGFET_HPNW8
XI6.X0 N_NET21_XI6.X0_D N_VDD_XI6.X0_PGD N_A_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW8
XI8.X0 N_Z_XI8.X0_D N_VDD_XI8.X0_PGD N_NET21_XI8.X0_CG N_VDD_XI8.X0_PGS
+ N_VSS_XI8.X0_S TIGFET_HPNW8
XI9.X0 N_Z_XI9.X0_D N_VSS_XI9.X0_PGD N_NET21_XI9.X0_CG N_VSS_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW8
*
x_PM_G3_OR2_N2_VSS N_VSS_XI7.X0_S N_VSS_XI5.X0_PGD N_VSS_XI6.X0_S N_VSS_XI8.X0_S
+ N_VSS_XI9.X0_PGD N_VSS_XI9.X0_PGS N_VSS_c_30_p N_VSS_c_4_p N_VSS_c_3_p
+ N_VSS_c_10_p N_VSS_c_53_p N_VSS_c_5_p N_VSS_c_8_p N_VSS_c_21_p N_VSS_c_28_p
+ N_VSS_c_15_p N_VSS_c_29_p N_VSS_c_6_p N_VSS_c_7_p VSS N_VSS_c_16_p
+ N_VSS_c_19_p N_VSS_c_17_p N_VSS_c_25_p N_VSS_c_18_p N_VSS_c_26_p Vss
+ PM_G3_OR2_N2_VSS
x_PM_G3_OR2_N2_VDD N_VDD_XI7.X0_PGD N_VDD_XI7.X0_PGS N_VDD_XI5.X0_S
+ N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI8.X0_PGD N_VDD_XI8.X0_PGS
+ N_VDD_XI9.X0_S N_VDD_c_72_n N_VDD_c_73_n N_VDD_c_114_p N_VDD_c_124_p
+ N_VDD_c_142_p N_VDD_c_74_n N_VDD_c_77_n N_VDD_c_79_n N_VDD_c_81_n N_VDD_c_82_n
+ N_VDD_c_88_n N_VDD_c_116_p N_VDD_c_89_n N_VDD_c_92_n N_VDD_c_96_n N_VDD_c_99_n
+ N_VDD_c_144_p N_VDD_c_104_n VDD N_VDD_c_107_n N_VDD_c_108_n N_VDD_c_109_n
+ N_VDD_c_117_p N_VDD_c_110_n N_VDD_c_112_n Vss PM_G3_OR2_N2_VDD
x_PM_G3_OR2_N2_B N_B_XI7.X0_CG N_B_XI5.X0_CG N_B_c_153_n N_B_c_165_p N_B_c_148_n
+ B N_B_c_157_n N_B_c_151_n Vss PM_G3_OR2_N2_B
x_PM_G3_OR2_N2_NET21 N_NET21_XI7.X0_D N_NET21_XI5.X0_D N_NET21_XI6.X0_D
+ N_NET21_XI8.X0_CG N_NET21_XI9.X0_CG N_NET21_c_169_n N_NET21_c_184_n
+ N_NET21_c_170_n N_NET21_c_172_n N_NET21_c_174_n N_NET21_c_179_n
+ N_NET21_c_194_n N_NET21_c_180_n Vss PM_G3_OR2_N2_NET21
x_PM_G3_OR2_N2_A N_A_XI5.X0_PGS N_A_XI6.X0_CG N_A_c_208_n N_A_c_211_n
+ N_A_c_213_n N_A_c_215_n A Vss PM_G3_OR2_N2_A
x_PM_G3_OR2_N2_Z N_Z_XI8.X0_D N_Z_XI9.X0_D N_Z_c_229_n Z N_Z_c_231_n Vss
+ PM_G3_OR2_N2_Z
cc_1 N_VSS_XI5.X0_PGD N_VDD_XI6.X0_PGD 0.00204282f
cc_2 N_VSS_XI9.X0_PGD N_VDD_XI8.X0_PGD 0.00196484f
cc_3 N_VSS_c_3_p N_VDD_c_72_n 0.00204282f
cc_4 N_VSS_c_4_p N_VDD_c_73_n 0.00196484f
cc_5 N_VSS_c_5_p N_VDD_c_74_n 0.00187494f
cc_6 N_VSS_c_6_p N_VDD_c_74_n 0.00677253f
cc_7 N_VSS_c_7_p N_VDD_c_74_n 0.00189302f
cc_8 N_VSS_c_8_p N_VDD_c_77_n 4.76491e-19
cc_9 N_VSS_c_6_p N_VDD_c_77_n 0.0033599f
cc_10 N_VSS_c_10_p N_VDD_c_79_n 3.44698e-19
cc_11 N_VSS_c_5_p N_VDD_c_79_n 9.72065e-19
cc_12 N_VSS_c_5_p N_VDD_c_81_n 4.54347e-19
cc_13 N_VSS_c_3_p N_VDD_c_82_n 3.66315e-19
cc_14 N_VSS_c_8_p N_VDD_c_82_n 0.00141228f
cc_15 N_VSS_c_15_p N_VDD_c_82_n 0.00114511f
cc_16 N_VSS_c_16_p N_VDD_c_82_n 0.00350144f
cc_17 N_VSS_c_17_p N_VDD_c_82_n 0.00435073f
cc_18 N_VSS_c_18_p N_VDD_c_82_n 7.74609e-19
cc_19 N_VSS_c_19_p N_VDD_c_88_n 0.00106851f
cc_20 N_VSS_c_8_p N_VDD_c_89_n 8.39054e-19
cc_21 N_VSS_c_21_p N_VDD_c_89_n 3.93845e-19
cc_22 N_VSS_c_15_p N_VDD_c_89_n 3.95933e-19
cc_23 N_VSS_c_21_p N_VDD_c_92_n 4.34701e-19
cc_24 N_VSS_c_17_p N_VDD_c_92_n 0.00137965f
cc_25 N_VSS_c_25_p N_VDD_c_92_n 0.00142692f
cc_26 N_VSS_c_26_p N_VDD_c_92_n 0.00107375f
cc_27 N_VSS_c_21_p N_VDD_c_96_n 3.91951e-19
cc_28 N_VSS_c_28_p N_VDD_c_96_n 8.45954e-19
cc_29 N_VSS_c_29_p N_VDD_c_96_n 3.99794e-19
cc_30 N_VSS_c_30_p N_VDD_c_99_n 4.1253e-19
cc_31 N_VSS_c_4_p N_VDD_c_99_n 3.9313e-19
cc_32 N_VSS_c_28_p N_VDD_c_99_n 0.00161703f
cc_33 N_VSS_c_29_p N_VDD_c_99_n 2.26455e-19
cc_34 N_VSS_c_25_p N_VDD_c_99_n 0.00609002f
cc_35 N_VSS_XI9.X0_PGS N_VDD_c_104_n 3.05236e-19
cc_36 N_VSS_c_28_p N_VDD_c_104_n 8.67538e-19
cc_37 N_VSS_c_29_p N_VDD_c_104_n 3.66936e-19
cc_38 N_VSS_c_6_p N_VDD_c_107_n 0.00116512f
cc_39 N_VSS_c_17_p N_VDD_c_108_n 9.95024e-19
cc_40 N_VSS_c_25_p N_VDD_c_109_n 9.97484e-19
cc_41 N_VSS_c_8_p N_VDD_c_110_n 3.44698e-19
cc_42 N_VSS_c_15_p N_VDD_c_110_n 6.36088e-19
cc_43 N_VSS_c_28_p N_VDD_c_112_n 3.48267e-19
cc_44 N_VSS_c_29_p N_VDD_c_112_n 6.489e-19
cc_45 N_VSS_c_8_p N_B_c_148_n 5.58916e-19
cc_46 N_VSS_c_15_p N_B_c_148_n 3.52408e-19
cc_47 N_VSS_c_6_p N_B_c_148_n 8.9847e-19
cc_48 N_VSS_c_8_p N_B_c_151_n 3.2351e-19
cc_49 N_VSS_c_15_p N_B_c_151_n 0.00119577f
cc_50 N_VSS_XI9.X0_PGD N_NET21_c_169_n 4.25712e-19
cc_51 N_VSS_c_10_p N_NET21_c_170_n 3.43419e-19
cc_52 N_VSS_c_5_p N_NET21_c_170_n 3.48267e-19
cc_53 N_VSS_c_53_p N_NET21_c_172_n 3.43419e-19
cc_54 N_VSS_c_21_p N_NET21_c_172_n 3.48267e-19
cc_55 N_VSS_c_10_p N_NET21_c_174_n 3.48267e-19
cc_56 N_VSS_c_53_p N_NET21_c_174_n 3.48267e-19
cc_57 N_VSS_c_5_p N_NET21_c_174_n 8.54909e-19
cc_58 N_VSS_c_21_p N_NET21_c_174_n 5.71987e-19
cc_59 N_VSS_c_6_p N_NET21_c_174_n 6.84771e-19
cc_60 N_VSS_c_25_p N_NET21_c_179_n 2.36784e-19
cc_61 N_VSS_c_21_p N_NET21_c_180_n 9.51297e-19
cc_62 N_VSS_c_6_p N_NET21_c_180_n 2.32409e-19
cc_63 N_VSS_c_17_p N_NET21_c_180_n 8.71002e-19
cc_64 N_VSS_XI5.X0_PGD N_A_c_208_n 9.55607e-19
cc_65 N_VSS_c_53_p N_Z_c_229_n 3.43419e-19
cc_66 N_VSS_c_21_p N_Z_c_229_n 3.48267e-19
cc_67 N_VSS_c_53_p N_Z_c_231_n 3.48267e-19
cc_68 N_VSS_c_21_p N_Z_c_231_n 7.85754e-19
cc_69 N_VSS_c_25_p N_Z_c_231_n 2.50289e-19
cc_70 N_VDD_c_114_p N_B_c_153_n 8.95172e-19
cc_71 N_VDD_c_74_n N_B_c_148_n 0.00268777f
cc_72 N_VDD_c_116_p N_B_c_148_n 5.04982e-19
cc_73 N_VDD_c_117_p N_B_c_148_n 3.55951e-19
cc_74 N_VDD_c_74_n N_B_c_157_n 5.06499e-19
cc_75 N_VDD_c_116_p N_B_c_157_n 3.47446e-19
cc_76 N_VDD_c_117_p N_B_c_157_n 2.75266e-19
cc_77 N_VDD_c_74_n N_B_c_151_n 3.66936e-19
cc_78 N_VDD_XI8.X0_PGD N_NET21_c_169_n 4.28909e-19
cc_79 N_VDD_c_112_n N_NET21_c_184_n 9.53212e-19
cc_80 N_VDD_c_124_p N_NET21_c_172_n 3.43419e-19
cc_81 N_VDD_c_81_n N_NET21_c_172_n 3.72199e-19
cc_82 N_VDD_c_82_n N_NET21_c_172_n 3.4118e-19
cc_83 N_VDD_c_124_p N_NET21_c_174_n 3.48267e-19
cc_84 N_VDD_c_74_n N_NET21_c_174_n 8.27149e-19
cc_85 N_VDD_c_81_n N_NET21_c_174_n 7.92786e-19
cc_86 N_VDD_c_82_n N_NET21_c_174_n 4.80596e-19
cc_87 N_VDD_c_96_n N_NET21_c_179_n 3.42685e-19
cc_88 N_VDD_c_112_n N_NET21_c_179_n 3.2351e-19
cc_89 N_VDD_c_112_n N_NET21_c_194_n 2.68747e-19
cc_90 N_VDD_XI7.X0_PGD N_A_c_208_n 5.1398e-19
cc_91 N_VDD_XI6.X0_PGD N_A_c_208_n 2.51476e-19
cc_92 N_VDD_XI7.X0_PGS N_A_c_211_n 6.75208e-19
cc_93 N_VDD_c_74_n N_A_c_211_n 4.39208e-19
cc_94 N_VDD_c_89_n N_A_c_213_n 3.47446e-19
cc_95 N_VDD_c_110_n N_A_c_213_n 0.00119807f
cc_96 N_VDD_c_89_n N_A_c_215_n 4.0116e-19
cc_97 N_VDD_c_110_n N_A_c_215_n 3.26762e-19
cc_98 N_VDD_c_142_p N_Z_c_229_n 3.43419e-19
cc_99 N_VDD_c_99_n N_Z_c_229_n 3.4118e-19
cc_100 N_VDD_c_144_p N_Z_c_229_n 3.72199e-19
cc_101 N_VDD_c_142_p N_Z_c_231_n 3.48267e-19
cc_102 N_VDD_c_99_n N_Z_c_231_n 4.63968e-19
cc_103 N_VDD_c_144_p N_Z_c_231_n 7.4527e-19
cc_104 N_B_c_148_n N_NET21_c_174_n 0.00749505f
cc_105 N_B_c_157_n N_NET21_c_174_n 0.0010409f
cc_106 N_B_c_151_n N_NET21_c_174_n 9.42705e-19
cc_107 N_B_c_148_n N_NET21_c_180_n 2.06853e-19
cc_108 N_B_c_165_p N_A_XI5.X0_PGS 5.00154e-19
cc_109 N_B_c_151_n N_A_XI5.X0_PGS 7.86826e-19
cc_110 N_B_c_157_n N_A_c_208_n 0.0015904f
cc_111 N_B_c_151_n N_A_c_213_n 7.50183e-19
cc_112 N_NET21_c_172_n N_A_c_208_n 4.45882e-19
cc_113 N_NET21_c_174_n N_A_c_208_n 8.51551e-19
cc_114 N_NET21_c_174_n N_A_c_213_n 0.00108501f
cc_115 N_NET21_c_179_n N_A_c_213_n 3.48267e-19
cc_116 N_NET21_c_194_n N_A_c_213_n 0.00171208f
cc_117 N_NET21_c_174_n N_A_c_215_n 0.0014331f
cc_118 N_NET21_c_179_n N_A_c_215_n 4.16154e-19
cc_119 N_NET21_c_180_n N_A_c_215_n 3.53251e-19
cc_120 N_NET21_c_169_n N_Z_c_229_n 6.55689e-19
*
.ends
*
*
.subckt OR2_HPNW8 A B Y VDD VSS
xgate (VSS VDD B A Y) G3_OR2_N2
.ends
*
* File: G4_XNOR2_N2.pex.netlist
* Created: Wed Mar 16 11:10:33 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XNOR2_N2_VDD 2 5 9 12 14 16 32 42 43 45 54 59 63 66 68 69 70 73 75
+ 76 79 81 85 89 91 93 98 99 100 103 109 114 Vss
c104 114 Vss 0.00451172f
c105 109 Vss 0.0046333f
c106 101 Vss 8.60971e-19
c107 100 Vss 2.39889e-19
c108 99 Vss 4.52364e-19
c109 98 Vss 0.00501239f
c110 93 Vss 0.00287584f
c111 91 Vss 0.0106993f
c112 89 Vss 0.00158164f
c113 85 Vss 4.92677e-19
c114 81 Vss 0.00450584f
c115 79 Vss 0.00110794f
c116 76 Vss 8.67986e-19
c117 75 Vss 0.00221168f
c118 73 Vss 0.00195091f
c119 70 Vss 8.63914e-19
c120 69 Vss 0.005504f
c121 68 Vss 0.00838153f
c122 66 Vss 0.00213842f
c123 63 Vss 0.00546856f
c124 59 Vss 0.00725053f
c125 54 Vss 0.00546856f
c126 45 Vss 1.15207e-19
c127 43 Vss 0.0351228f
c128 42 Vss 0.100955f
c129 33 Vss 0.035919f
c130 32 Vss 0.100953f
c131 14 Vss 0.00143442f
c132 9 Vss 0.266831f
c133 5 Vss 0.270069f
r134 98 103 0.326018
r135 97 98 4.58464
r136 93 97 0.655813
r137 93 95 1.82344
r138 92 101 0.494161
r139 91 103 0.326018
r140 91 92 13.0037
r141 87 101 0.128424
r142 87 89 5.2515
r143 85 114 1.16709
r144 83 85 2.16729
r145 82 100 0.494161
r146 81 101 0.494161
r147 81 82 7.46046
r148 79 109 1.16709
r149 77 100 0.128424
r150 77 79 2.16729
r151 75 100 0.494161
r152 75 76 4.37625
r153 71 99 0.0828784
r154 71 73 1.82344
r155 69 83 0.652036
r156 69 70 10.1279
r157 68 76 0.652036
r158 67 99 0.551426
r159 67 68 14.7125
r160 66 99 0.551426
r161 65 70 0.652036
r162 65 66 4.58464
r163 63 95 1.16709
r164 59 89 1.16709
r165 54 73 1.16709
r166 45 114 0.0476429
r167 43 45 1.45875
r168 42 46 0.652036
r169 42 45 1.45875
r170 39 43 0.652036
r171 35 109 0.0476429
r172 33 35 1.45875
r173 32 36 0.652036
r174 32 35 1.45875
r175 29 33 0.652036
r176 16 63 0.185659
r177 14 59 0.185659
r178 12 59 0.185659
r179 9 46 3.8511
r180 9 39 3.8511
r181 5 36 3.8511
r182 5 29 3.8511
r183 2 54 0.185659
.ends

.subckt PM_G4_XNOR2_N2_VSS 3 6 8 11 14 16 32 33 42 43 54 59 63 66 71 76 81 87 96
+ 101 114 116 117 118 123 124 129 137 142 143 144 146 Vss
c87 144 Vss 3.75522e-19
c88 143 Vss 4.28045e-19
c89 142 Vss 0.00380395f
c90 137 Vss 0.00119929f
c91 129 Vss 0.0129925f
c92 124 Vss 8.20954e-19
c93 123 Vss 0.00416713f
c94 118 Vss 8.42922e-19
c95 117 Vss 0.00171404f
c96 116 Vss 0.00154361f
c97 114 Vss 0.00516329f
c98 101 Vss 0.00400427f
c99 96 Vss 0.00412244f
c100 87 Vss 1.41859e-19
c101 81 Vss 0.00270839f
c102 76 Vss 8.07404e-19
c103 71 Vss 0.00125472f
c104 66 Vss 0.00178947f
c105 63 Vss 0.00389308f
c106 59 Vss 0.00728678f
c107 54 Vss 0.0039211f
c108 43 Vss 0.0342891f
c109 42 Vss 0.100066f
c110 35 Vss 1.95386e-19
c111 33 Vss 0.0350852f
c112 32 Vss 0.0990713f
c113 14 Vss 0.00143442f
c114 11 Vss 0.269838f
c115 3 Vss 0.266926f
r116 142 146 0.349767
r117 141 142 4.58464
r118 137 146 0.306046
r119 130 144 0.494161
r120 129 141 0.652036
r121 125 144 0.128424
r122 123 133 0.652036
r123 123 124 10.1279
r124 119 143 0.0828784
r125 117 144 0.494161
r126 117 118 4.37625
r127 116 124 0.652036
r128 115 143 0.551426
r129 115 116 4.58464
r130 114 143 0.551426
r131 113 118 0.652036
r132 113 114 14.7125
r133 87 137 1.82344
r134 81 129 13.5872
r135 81 130 8.04396
r136 81 84 5.79332
r137 76 101 1.16709
r138 76 133 2.16729
r139 71 96 1.16709
r140 71 125 2.16729
r141 66 119 1.82344
r142 63 87 1.16709
r143 59 84 1.16709
r144 54 66 1.16709
r145 45 101 0.0476429
r146 43 45 1.45875
r147 42 46 0.652036
r148 42 45 1.45875
r149 39 43 0.652036
r150 35 96 0.0476429
r151 33 35 1.45875
r152 32 36 0.652036
r153 32 35 1.45875
r154 29 33 0.652036
r155 16 63 0.185659
r156 14 59 0.185659
r157 11 46 3.8511
r158 11 39 3.8511
r159 8 59 0.185659
r160 6 54 0.185659
r161 3 36 3.8511
r162 3 29 3.8511
.ends

.subckt PM_G4_XNOR2_N2_A 2 4 7 10 21 24 28 39 48 53 56 61 66 71 76 84 Vss
c57 84 Vss 4.74028e-19
c58 76 Vss 8.09766e-19
c59 71 Vss 0.00526551f
c60 66 Vss 0.00379683f
c61 61 Vss 0.00265207f
c62 56 Vss 0.0049943f
c63 53 Vss 8.5599e-19
c64 48 Vss 0.126052f
c65 43 Vss 0.0296526f
c66 39 Vss 1.95944e-19
c67 28 Vss 0.152877f
c68 24 Vss 1.05421e-19
c69 21 Vss 0.169632f
c70 18 Vss 0.12596f
c71 16 Vss 0.0247918f
c72 10 Vss 0.121972f
c73 7 Vss 0.324361f
c74 4 Vss 0.138512f
r75 80 84 0.652036
r76 61 76 1.16709
r77 61 84 5.20982
r78 56 71 1.16709
r79 56 80 9.54439
r80 53 66 1.16709
r81 47 71 0.0238214
r82 47 48 2.334
r83 44 47 2.20433
r84 39 76 0.404964
r85 33 48 0.00605528
r86 31 44 0.00605528
r87 29 43 0.494161
r88 28 30 0.652036
r89 28 29 4.84305
r90 25 43 0.128424
r91 24 66 0.0476429
r92 22 24 0.326018
r93 22 24 0.1167
r94 21 43 0.494161
r95 21 24 6.7686
r96 18 66 0.357321
r97 16 24 0.326018
r98 16 18 0.40845
r99 10 39 3.32595
r100 7 33 3.8511
r101 7 31 3.8511
r102 7 30 3.8511
r103 4 25 3.8511
r104 2 18 3.44265
.ends

.subckt PM_G4_XNOR2_N2_NET1 2 4 7 10 30 31 35 41 44 49 58 66 Vss
c34 66 Vss 2.19199e-19
c35 58 Vss 0.0058571f
c36 49 Vss 0.00612925f
c37 44 Vss 0.00128347f
c38 41 Vss 0.00534332f
c39 35 Vss 0.103384f
c40 31 Vss 0.12896f
c41 30 Vss 1.02017e-19
c42 10 Vss 0.236304f
c43 7 Vss 0.381296f
c44 4 Vss 0.00143442f
r45 62 66 0.652036
r46 49 58 1.16709
r47 49 66 13.8373
r48 44 62 2.50071
r49 41 44 1.16709
r50 33 35 1.70187
r51 30 58 0.0238214
r52 30 31 2.20433
r53 27 30 2.334
r54 25 35 0.17282
r55 24 31 0.00605528
r56 21 33 0.17282
r57 18 27 0.00605528
r58 10 21 7.06035
r59 7 25 5.7183
r60 7 24 3.8511
r61 7 18 3.8511
r62 4 41 0.185659
r63 2 41 0.185659
.ends

.subckt PM_G4_XNOR2_N2_NET3 2 4 6 9 21 22 33 39 42 47 56 74 Vss
c49 74 Vss 3.4517e-19
c50 56 Vss 0.0039047f
c51 47 Vss 0.00714759f
c52 42 Vss 0.00198779f
c53 39 Vss 0.00534332f
c54 33 Vss 0.12548f
c55 22 Vss 0.0340569f
c56 21 Vss 0.175814f
c57 9 Vss 0.464757f
c58 6 Vss 0.145805f
c59 4 Vss 0.00143442f
r60 70 74 0.655813
r61 47 56 1.16709
r62 47 74 12.0712
r63 42 70 2.41736
r64 39 42 1.16709
r65 32 56 0.0238214
r66 32 33 2.26917
r67 29 32 2.26917
r68 26 33 0.00605528
r69 24 29 0.00605528
r70 21 23 0.652036
r71 21 22 4.84305
r72 18 22 0.652036
r73 9 26 3.8511
r74 9 24 3.8511
r75 9 23 8.7525
r76 6 18 4.25955
r77 4 39 0.185659
r78 2 39 0.185659
.ends

.subckt PM_G4_XNOR2_N2_B 2 4 7 10 19 20 28 31 33 37 38 48 52 58 61 Vss
c36 61 Vss 0.0281739f
c37 58 Vss 0.00110612f
c38 52 Vss 0.136411f
c39 48 Vss 0.0595342f
c40 38 Vss 0.0333783f
c41 37 Vss 0.090268f
c42 33 Vss 0.0442143f
c43 31 Vss 9.80304e-20
c44 28 Vss 0.0899896f
c45 20 Vss 0.0348277f
c46 19 Vss 0.169632f
c47 10 Vss 0.209756f
c48 7 Vss 0.322768f
c49 4 Vss 0.125964f
c50 2 Vss 0.138383f
r51 55 61 1.16709
r52 55 58 0.0729375
r53 50 52 4.53833
r54 47 48 1.167
r55 42 52 0.00605528
r56 37 39 0.652036
r57 37 38 2.04225
r58 35 48 0.0685365
r59 34 50 0.00605528
r60 33 38 0.652036
r61 32 47 0.0685365
r62 32 33 1.69215
r63 31 61 0.181909
r64 29 61 0.494161
r65 29 31 0.1167
r66 28 47 0.5835
r67 28 31 3.55935
r68 23 61 0.128424
r69 23 61 0.40845
r70 22 61 0.181909
r71 20 22 6.7686
r72 19 61 0.494161
r73 19 22 0.1167
r74 16 20 0.652036
r75 10 39 6.3018
r76 7 42 3.8511
r77 7 35 3.8511
r78 7 34 3.8511
r79 4 61 3.44265
r80 2 16 3.8511
.ends

.subckt PM_G4_XNOR2_N2_Z 2 4 6 8 23 27 30 33 Vss
c29 30 Vss 0.00338645f
c30 27 Vss 0.0063256f
c31 23 Vss 0.00620875f
c32 8 Vss 0.00143442f
c33 6 Vss 0.00143442f
r34 33 35 4.668
r35 30 33 5.45989
r36 27 35 1.16709
r37 23 30 1.16709
r38 8 27 0.185659
r39 6 23 0.185659
r40 4 27 0.185659
r41 2 23 0.185659
.ends

.subckt G4_XNOR2_N2  VDD VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI16.X0 N_NET1_XI16.X0_D N_VSS_XI16.X0_PGD N_B_XI16.X0_CG N_VSS_XI16.X0_PGD
+ N_VDD_XI16.X0_S TIGFET_HPNW8
XI12.X0 N_NET3_XI12.X0_D N_VDD_XI12.X0_PGD N_A_XI12.X0_CG N_VDD_XI12.X0_PGD
+ N_VSS_XI12.X0_S TIGFET_HPNW8
XI18.X0 N_NET1_XI18.X0_D N_VDD_XI18.X0_PGD N_B_XI18.X0_CG N_VDD_XI18.X0_PGD
+ N_VSS_XI18.X0_S TIGFET_HPNW8
XI13.X0 N_NET3_XI13.X0_D N_VSS_XI13.X0_PGD N_A_XI13.X0_CG N_VSS_XI13.X0_PGD
+ N_VDD_XI13.X0_S TIGFET_HPNW8
XI17.X0 N_Z_XI17.X0_D N_B_XI17.X0_PGD N_NET3_XI17.X0_CG N_B_XI17.X0_PGD
+ N_VSS_XI17.X0_S TIGFET_HPNW8
XI14.X0 N_Z_XI14.X0_D N_A_XI14.X0_PGD N_B_XI14.X0_CG N_A_XI14.X0_PGD
+ N_VDD_XI14.X0_S TIGFET_HPNW8
XI19.X0 N_Z_XI19.X0_D N_NET1_XI19.X0_PGD N_A_XI19.X0_CG N_NET1_XI19.X0_PGD
+ N_VSS_XI19.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_NET3_XI15.X0_PGD N_NET1_XI15.X0_CG N_NET3_XI15.X0_PGD
+ N_VDD_XI15.X0_S TIGFET_HPNW8
*
x_PM_G4_XNOR2_N2_VDD N_VDD_XI16.X0_S N_VDD_XI12.X0_PGD N_VDD_XI18.X0_PGD
+ N_VDD_XI13.X0_S N_VDD_XI14.X0_S N_VDD_XI15.X0_S N_VDD_c_9_p N_VDD_c_23_p
+ N_VDD_c_5_p N_VDD_c_89_p N_VDD_c_65_p N_VDD_c_11_p N_VDD_c_96_p N_VDD_c_7_p
+ N_VDD_c_12_p N_VDD_c_6_p N_VDD_c_40_p N_VDD_c_13_p N_VDD_c_14_p N_VDD_c_44_p
+ N_VDD_c_19_p N_VDD_c_10_p N_VDD_c_17_p N_VDD_c_4_p N_VDD_c_54_p N_VDD_c_27_p
+ N_VDD_c_72_p N_VDD_c_37_p N_VDD_c_43_p VDD N_VDD_c_22_p N_VDD_c_18_p Vss
+ PM_G4_XNOR2_N2_VDD
x_PM_G4_XNOR2_N2_VSS N_VSS_XI16.X0_PGD N_VSS_XI12.X0_S N_VSS_XI18.X0_S
+ N_VSS_XI13.X0_PGD N_VSS_XI17.X0_S N_VSS_XI19.X0_S N_VSS_c_109_n N_VSS_c_111_n
+ N_VSS_c_157_p N_VSS_c_113_n N_VSS_c_173_p N_VSS_c_115_n N_VSS_c_185_p
+ N_VSS_c_116_n N_VSS_c_119_n N_VSS_c_123_n N_VSS_c_127_n N_VSS_c_131_n
+ N_VSS_c_132_n N_VSS_c_136_n N_VSS_c_139_n N_VSS_c_142_n N_VSS_c_143_n
+ N_VSS_c_144_n N_VSS_c_145_n N_VSS_c_148_n N_VSS_c_149_n N_VSS_c_150_n
+ N_VSS_c_169_p N_VSS_c_151_n N_VSS_c_152_n VSS Vss PM_G4_XNOR2_N2_VSS
x_PM_G4_XNOR2_N2_A N_A_XI12.X0_CG N_A_XI13.X0_CG N_A_XI14.X0_PGD N_A_XI19.X0_CG
+ N_A_c_193_n N_A_c_195_n N_A_c_196_n N_A_c_220_p N_A_c_197_n A N_A_c_201_n
+ N_A_c_221_p N_A_c_203_n N_A_c_206_n N_A_c_219_p N_A_c_217_n Vss
+ PM_G4_XNOR2_N2_A
x_PM_G4_XNOR2_N2_NET1 N_NET1_XI16.X0_D N_NET1_XI18.X0_D N_NET1_XI19.X0_PGD
+ N_NET1_XI15.X0_CG N_NET1_c_268_n N_NET1_c_281_p N_NET1_c_274_p N_NET1_c_249_n
+ N_NET1_c_252_n N_NET1_c_255_n N_NET1_c_271_n N_NET1_c_263_n Vss
+ PM_G4_XNOR2_N2_NET1
x_PM_G4_XNOR2_N2_NET3 N_NET3_XI12.X0_D N_NET3_XI13.X0_D N_NET3_XI17.X0_CG
+ N_NET3_XI15.X0_PGD N_NET3_c_306_n N_NET3_c_323_p N_NET3_c_284_n N_NET3_c_285_n
+ N_NET3_c_286_n N_NET3_c_289_n N_NET3_c_292_n N_NET3_c_294_n Vss
+ PM_G4_XNOR2_N2_NET3
x_PM_G4_XNOR2_N2_B N_B_XI16.X0_CG N_B_XI18.X0_CG N_B_XI17.X0_PGD N_B_XI14.X0_CG
+ N_B_c_334_n N_B_c_349_n N_B_c_336_n N_B_c_337_n N_B_c_361_n N_B_c_357_n
+ N_B_c_351_n N_B_c_365_n N_B_c_338_n B N_B_c_341_n Vss PM_G4_XNOR2_N2_B
x_PM_G4_XNOR2_N2_Z N_Z_XI17.X0_D N_Z_XI14.X0_D N_Z_XI19.X0_D N_Z_XI15.X0_D
+ N_Z_c_378_n N_Z_c_368_n N_Z_c_373_n Z Vss PM_G4_XNOR2_N2_Z
cc_1 N_VDD_XI12.X0_PGD N_VSS_XI16.X0_PGD 2.89249e-19
cc_2 N_VDD_XI18.X0_PGD N_VSS_XI16.X0_PGD 0.00196286f
cc_3 N_VDD_XI12.X0_PGD N_VSS_XI13.X0_PGD 0.0019593f
cc_4 N_VDD_c_4_p N_VSS_XI13.X0_PGD 2.22629e-19
cc_5 N_VDD_c_5_p N_VSS_c_109_n 0.00196286f
cc_6 N_VDD_c_6_p N_VSS_c_109_n 3.9313e-19
cc_7 N_VDD_c_7_p N_VSS_c_111_n 2.76462e-19
cc_8 N_VDD_c_6_p N_VSS_c_111_n 3.9313e-19
cc_9 N_VDD_c_9_p N_VSS_c_113_n 0.0019593f
cc_10 N_VDD_c_10_p N_VSS_c_113_n 3.9313e-19
cc_11 N_VDD_c_11_p N_VSS_c_115_n 3.13688e-19
cc_12 N_VDD_c_12_p N_VSS_c_116_n 0.00187494f
cc_13 N_VDD_c_13_p N_VSS_c_116_n 5.06564e-19
cc_14 N_VDD_c_14_p N_VSS_c_116_n 4.5625e-19
cc_15 N_VDD_c_7_p N_VSS_c_119_n 4.35319e-19
cc_16 N_VDD_c_6_p N_VSS_c_119_n 0.00141228f
cc_17 N_VDD_c_17_p N_VSS_c_119_n 8.69067e-19
cc_18 N_VDD_c_18_p N_VSS_c_119_n 3.48267e-19
cc_19 N_VDD_c_19_p N_VSS_c_123_n 9.53862e-19
cc_20 N_VDD_c_10_p N_VSS_c_123_n 0.00161703f
cc_21 N_VDD_c_4_p N_VSS_c_123_n 0.00227772f
cc_22 N_VDD_c_22_p N_VSS_c_123_n 3.48267e-19
cc_23 N_VDD_c_23_p N_VSS_c_127_n 2.38046e-19
cc_24 N_VDD_c_6_p N_VSS_c_127_n 0.00534412f
cc_25 N_VDD_c_4_p N_VSS_c_127_n 3.34043e-19
cc_26 N_VDD_c_18_p N_VSS_c_127_n 9.58524e-19
cc_27 N_VDD_c_27_p N_VSS_c_131_n 2.11881e-19
cc_28 N_VDD_c_7_p N_VSS_c_132_n 3.66936e-19
cc_29 N_VDD_c_6_p N_VSS_c_132_n 0.00114511f
cc_30 N_VDD_c_17_p N_VSS_c_132_n 3.99794e-19
cc_31 N_VDD_c_18_p N_VSS_c_132_n 6.489e-19
cc_32 N_VDD_c_10_p N_VSS_c_136_n 2.26455e-19
cc_33 N_VDD_c_4_p N_VSS_c_136_n 9.55322e-19
cc_34 N_VDD_c_22_p N_VSS_c_136_n 6.46219e-19
cc_35 N_VDD_c_7_p N_VSS_c_139_n 0.00309754f
cc_36 N_VDD_c_12_p N_VSS_c_139_n 0.00766101f
cc_37 N_VDD_c_37_p N_VSS_c_139_n 0.0010706f
cc_38 N_VDD_c_12_p N_VSS_c_142_n 0.0033176f
cc_39 N_VDD_c_6_p N_VSS_c_143_n 0.00345383f
cc_40 N_VDD_c_40_p N_VSS_c_144_n 0.00107685f
cc_41 N_VDD_c_14_p N_VSS_c_145_n 0.0035394f
cc_42 N_VDD_c_10_p N_VSS_c_145_n 0.00604286f
cc_43 N_VDD_c_43_p N_VSS_c_145_n 0.00103916f
cc_44 N_VDD_c_44_p N_VSS_c_148_n 0.0010609f
cc_45 N_VDD_c_6_p N_VSS_c_149_n 0.00459995f
cc_46 N_VDD_c_27_p N_VSS_c_150_n 0.00107435f
cc_47 N_VDD_c_12_p N_VSS_c_151_n 9.16632e-19
cc_48 N_VDD_c_6_p N_VSS_c_152_n 7.74609e-19
cc_49 N_VDD_c_4_p N_A_XI14.X0_PGD 2.06119e-19
cc_50 N_VDD_XI12.X0_PGD N_A_c_193_n 4.07423e-19
cc_51 N_VDD_XI18.X0_PGD N_A_c_193_n 2.2186e-19
cc_52 N_VDD_c_22_p N_A_c_195_n 9.45508e-19
cc_53 N_VDD_XI18.X0_PGD N_A_c_196_n 2.2186e-19
cc_54 N_VDD_c_54_p N_A_c_197_n 6.28504e-19
cc_55 N_VDD_c_12_p A 5.04211e-19
cc_56 N_VDD_c_19_p A 4.35492e-19
cc_57 N_VDD_c_22_p A 3.2351e-19
cc_58 N_VDD_c_4_p N_A_c_201_n 0.00256103f
cc_59 N_VDD_c_54_p N_A_c_201_n 0.00191796f
cc_60 N_VDD_c_12_p N_A_c_203_n 6.26183e-19
cc_61 N_VDD_c_19_p N_A_c_203_n 3.43988e-19
cc_62 N_VDD_c_22_p N_A_c_203_n 2.68747e-19
cc_63 N_VDD_c_4_p N_A_c_206_n 9.84209e-19
cc_64 N_VDD_c_54_p N_A_c_206_n 2.68554e-19
cc_65 N_VDD_c_65_p N_NET1_c_249_n 3.43419e-19
cc_66 N_VDD_c_6_p N_NET1_c_249_n 3.4118e-19
cc_67 N_VDD_c_13_p N_NET1_c_249_n 3.72199e-19
cc_68 N_VDD_c_65_p N_NET1_c_252_n 3.48267e-19
cc_69 N_VDD_c_6_p N_NET1_c_252_n 3.98099e-19
cc_70 N_VDD_c_13_p N_NET1_c_252_n 5.226e-19
cc_71 N_VDD_c_17_p N_NET1_c_255_n 0.00115819f
cc_72 N_VDD_c_72_p N_NET3_XI15.X0_PGD 2.91063e-19
cc_73 N_VDD_c_54_p N_NET3_c_284_n 8.60495e-19
cc_74 N_VDD_c_11_p N_NET3_c_285_n 3.43419e-19
cc_75 N_VDD_c_11_p N_NET3_c_286_n 3.48267e-19
cc_76 N_VDD_c_10_p N_NET3_c_286_n 4.34701e-19
cc_77 N_VDD_c_4_p N_NET3_c_286_n 0.00100809f
cc_78 N_VDD_c_4_p N_NET3_c_289_n 0.00119634f
cc_79 N_VDD_c_54_p N_NET3_c_289_n 0.00298078f
cc_80 N_VDD_c_72_p N_NET3_c_289_n 7.77543e-19
cc_81 N_VDD_c_54_p N_NET3_c_292_n 0.00118178f
cc_82 N_VDD_c_72_p N_NET3_c_292_n 3.66936e-19
cc_83 N_VDD_c_19_p N_NET3_c_294_n 2.94103e-19
cc_84 N_VDD_c_12_p N_B_XI16.X0_CG 2.61808e-19
cc_85 N_VDD_XI18.X0_PGD N_B_XI17.X0_PGD 0.00190378f
cc_86 N_VDD_XI12.X0_PGD N_B_c_334_n 2.2186e-19
cc_87 N_VDD_XI18.X0_PGD N_B_c_334_n 4.07423e-19
cc_88 N_VDD_XI18.X0_PGD N_B_c_336_n 4.08222e-19
cc_89 N_VDD_c_89_p N_B_c_337_n 9.08628e-19
cc_90 N_VDD_c_23_p N_B_c_338_n 0.00168656f
cc_91 N_VDD_c_17_p B 3.02102e-19
cc_92 N_VDD_c_18_p B 3.2351e-19
cc_93 N_VDD_c_17_p N_B_c_341_n 3.36818e-19
cc_94 N_VDD_c_18_p N_B_c_341_n 2.68747e-19
cc_95 N_VDD_c_11_p N_Z_c_368_n 3.43419e-19
cc_96 N_VDD_c_96_p N_Z_c_368_n 3.43419e-19
cc_97 N_VDD_c_4_p N_Z_c_368_n 3.48267e-19
cc_98 N_VDD_c_54_p N_Z_c_368_n 3.4118e-19
cc_99 N_VDD_c_27_p N_Z_c_368_n 3.72199e-19
cc_100 N_VDD_c_11_p N_Z_c_373_n 3.48267e-19
cc_101 N_VDD_c_96_p N_Z_c_373_n 3.48267e-19
cc_102 N_VDD_c_4_p N_Z_c_373_n 4.85404e-19
cc_103 N_VDD_c_54_p N_Z_c_373_n 5.96492e-19
cc_104 N_VDD_c_27_p N_Z_c_373_n 8.21216e-19
cc_105 N_VSS_XI13.X0_PGD N_A_XI14.X0_PGD 0.00164979f
cc_106 N_VSS_XI16.X0_PGD N_A_c_193_n 2.2186e-19
cc_107 N_VSS_XI13.X0_PGD N_A_c_193_n 4.04227e-19
cc_108 N_VSS_XI13.X0_PGD N_A_c_196_n 4.08222e-19
cc_109 N_VSS_c_157_p N_A_c_197_n 0.00164979f
cc_110 N_VSS_c_123_n N_A_c_201_n 3.87149e-19
cc_111 N_VSS_c_139_n N_A_c_201_n 4.99859e-19
cc_112 N_VSS_c_132_n N_A_c_203_n 2.38312e-19
cc_113 N_VSS_c_136_n N_A_c_206_n 6.52904e-19
cc_114 N_VSS_c_149_n N_A_c_217_n 6.07247e-19
cc_115 N_VSS_c_115_n N_NET1_c_249_n 3.43419e-19
cc_116 N_VSS_c_127_n N_NET1_c_249_n 3.48267e-19
cc_117 N_VSS_c_115_n N_NET1_c_252_n 3.48267e-19
cc_118 N_VSS_c_127_n N_NET1_c_252_n 0.00138658f
cc_119 N_VSS_c_127_n N_NET1_c_255_n 0.00157945f
cc_120 N_VSS_c_149_n N_NET1_c_255_n 0.0182344f
cc_121 N_VSS_c_169_p N_NET1_c_255_n 0.0011475f
cc_122 N_VSS_c_119_n N_NET1_c_263_n 0.00193107f
cc_123 N_VSS_c_139_n N_NET1_c_263_n 0.00107322f
cc_124 N_VSS_c_149_n N_NET1_c_263_n 0.00164616f
cc_125 N_VSS_c_173_p N_NET3_c_285_n 3.43419e-19
cc_126 N_VSS_c_173_p N_NET3_c_286_n 3.48267e-19
cc_127 N_VSS_c_116_n N_NET3_c_286_n 0.0011211f
cc_128 N_VSS_c_142_n N_NET3_c_286_n 4.15771e-19
cc_129 N_VSS_c_145_n N_NET3_c_286_n 2.79692e-19
cc_130 N_VSS_c_123_n N_NET3_c_289_n 0.00136387f
cc_131 N_VSS_c_145_n N_NET3_c_294_n 4.73555e-19
cc_132 N_VSS_XI16.X0_PGD N_B_c_334_n 4.04227e-19
cc_133 N_VSS_XI13.X0_PGD N_B_c_334_n 2.2186e-19
cc_134 N_VSS_XI13.X0_PGD N_B_c_336_n 2.2186e-19
cc_135 N_VSS_c_127_n N_B_c_338_n 2.49315e-19
cc_136 N_VSS_c_115_n N_Z_c_378_n 3.43419e-19
cc_137 N_VSS_c_185_p N_Z_c_378_n 3.43419e-19
cc_138 N_VSS_c_127_n N_Z_c_378_n 3.48267e-19
cc_139 N_VSS_c_131_n N_Z_c_378_n 3.48267e-19
cc_140 N_VSS_c_115_n N_Z_c_373_n 3.48267e-19
cc_141 N_VSS_c_185_p N_Z_c_373_n 3.48267e-19
cc_142 N_VSS_c_127_n N_Z_c_373_n 8.69457e-19
cc_143 N_VSS_c_131_n N_Z_c_373_n 5.71987e-19
cc_144 N_A_XI19.X0_CG N_NET1_XI19.X0_PGD 5.00154e-19
cc_145 N_A_c_219_p N_NET1_XI19.X0_PGD 0.00253213f
cc_146 N_A_c_220_p N_NET1_c_268_n 9.11431e-19
cc_147 N_A_c_221_p N_NET1_c_255_n 0.00300988f
cc_148 N_A_c_217_n N_NET1_c_255_n 8.60245e-19
cc_149 N_A_c_221_p N_NET1_c_271_n 3.14782e-19
cc_150 N_A_c_219_p N_NET1_c_271_n 2.68747e-19
cc_151 N_A_c_219_p N_NET3_XI17.X0_CG 2.16281e-19
cc_152 N_A_XI14.X0_PGD N_NET3_XI15.X0_PGD 0.00174198f
cc_153 N_A_c_196_n N_NET3_XI15.X0_PGD 3.14428e-19
cc_154 N_A_c_219_p N_NET3_XI15.X0_PGD 4.34237e-19
cc_155 N_A_XI14.X0_PGD N_NET3_c_306_n 4.63684e-19
cc_156 N_A_c_197_n N_NET3_c_284_n 0.00174198f
cc_157 N_A_c_193_n N_NET3_c_285_n 6.32063e-19
cc_158 N_A_c_201_n N_NET3_c_286_n 9.99037e-19
cc_159 N_A_c_201_n N_NET3_c_289_n 0.00251926f
cc_160 N_A_c_221_p N_NET3_c_289_n 0.00147102f
cc_161 N_A_c_206_n N_NET3_c_289_n 3.44698e-19
cc_162 N_A_c_220_p N_NET3_c_292_n 4.02896e-19
cc_163 N_A_c_201_n N_NET3_c_292_n 3.44698e-19
cc_164 N_A_c_206_n N_NET3_c_292_n 6.70706e-19
cc_165 N_A_c_196_n N_B_XI14.X0_CG 0.003858f
cc_166 N_A_c_193_n N_B_c_334_n 0.00500727f
cc_167 N_A_c_203_n N_B_c_349_n 6.36314e-19
cc_168 N_A_c_196_n N_B_c_336_n 0.00268264f
cc_169 N_A_c_196_n N_B_c_351_n 0.00354125f
cc_170 N_A_c_217_n B 2.16641e-19
cc_171 N_A_c_193_n N_B_c_341_n 0.00152783f
cc_172 N_A_c_201_n N_Z_c_373_n 0.00406991f
cc_173 N_A_c_221_p N_Z_c_373_n 0.00267623f
cc_174 N_A_c_219_p N_Z_c_373_n 0.00100289f
cc_175 N_NET1_XI19.X0_PGD N_NET3_XI17.X0_CG 3.24817e-19
cc_176 N_NET1_c_274_p N_NET3_XI15.X0_PGD 0.00863799f
cc_177 N_NET1_XI19.X0_PGD N_NET3_c_306_n 0.00333245f
cc_178 N_NET1_c_249_n N_NET3_c_285_n 2.31842e-19
cc_179 N_NET1_XI19.X0_PGD N_B_XI17.X0_PGD 0.00216194f
cc_180 N_NET1_XI15.X0_CG N_B_XI14.X0_CG 2.72501e-19
cc_181 N_NET1_c_249_n N_B_c_334_n 6.32063e-19
cc_182 N_NET1_c_274_p N_B_c_357_n 2.72501e-19
cc_183 N_NET1_c_281_p N_B_c_338_n 0.00193608f
cc_184 N_NET1_c_255_n N_Z_c_373_n 3.07539e-19
cc_185 N_NET3_XI17.X0_CG N_B_XI17.X0_PGD 0.00201028f
cc_186 N_NET3_c_306_n N_B_XI17.X0_PGD 0.00163252f
cc_187 N_NET3_XI15.X0_PGD N_B_c_361_n 3.23792e-19
cc_188 N_NET3_c_323_p N_B_c_361_n 5.75886e-19
cc_189 N_NET3_XI15.X0_PGD N_B_c_357_n 0.00310335f
cc_190 N_NET3_c_323_p N_B_c_357_n 0.00192667f
cc_191 N_NET3_c_323_p N_B_c_365_n 0.00201028f
cc_192 N_NET3_c_306_n N_Z_c_378_n 6.54859e-19
cc_193 N_NET3_c_306_n N_Z_c_368_n 2.54846e-19
cc_194 N_NET3_XI15.X0_PGD N_Z_c_373_n 0.00129454f
cc_195 N_NET3_c_306_n N_Z_c_373_n 2.46041e-19
cc_196 N_NET3_c_289_n N_Z_c_373_n 2.36895e-19
cc_197 N_B_c_357_n N_Z_c_373_n 9.47639e-19
cc_198 B N_Z_c_373_n 2.02757e-19
*
.ends
*
*
.subckt XNOR2_HPNW8 A B Y VDD VSS
xgate (VDD VSS A B Y) G4_XNOR2_N2
.ends
*
* File: G5_XNOR3_N2.pex.netlist
* Created: Mon Mar 28 15:31:24 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XNOR3_N2_VDD 2 3 5 8 10 11 29 30 41 42 44 53 54 65 69 74 83 85 86
+ 87 90 92 96 99 102 104 108 110 114 118 120 122 124 125 131 140 145 Vss
c116 145 Vss 0.00470693f
c117 140 Vss 0.00487376f
c118 131 Vss 0.00472091f
c119 125 Vss 2.39889e-19
c120 124 Vss 4.91772e-19
c121 123 Vss 5.21614e-19
c122 120 Vss 4.52364e-19
c123 118 Vss 0.00162316f
c124 114 Vss 4.81041e-19
c125 110 Vss 0.00631991f
c126 108 Vss 9.42823e-19
c127 104 Vss 0.00578311f
c128 102 Vss 0.00174133f
c129 99 Vss 0.00271006f
c130 96 Vss 0.00486611f
c131 92 Vss 0.00657264f
c132 90 Vss 0.00151669f
c133 87 Vss 8.67714e-19
c134 86 Vss 0.0090076f
c135 85 Vss 0.0105886f
c136 83 Vss 0.00212071f
c137 74 Vss 0.00377995f
c138 69 Vss 0.0039448f
c139 65 Vss 0.00373195f
c140 54 Vss 0.035607f
c141 53 Vss 0.100823f
c142 44 Vss 8.7772e-20
c143 42 Vss 0.0356105f
c144 41 Vss 0.101295f
c145 30 Vss 0.0346327f
c146 29 Vss 0.0990915f
c147 11 Vss 0.269218f
c148 5 Vss 0.27009f
c149 3 Vss 0.232895f
r150 116 118 5.2515
r151 114 145 1.16709
r152 112 114 2.16729
r153 111 125 0.494161
r154 110 116 0.652036
r155 110 111 7.46046
r156 108 140 1.16709
r157 106 125 0.128424
r158 106 108 2.16729
r159 105 124 0.494161
r160 104 112 0.652036
r161 104 105 10.3363
r162 100 123 0.0828784
r163 100 102 2.00578
r164 99 124 0.128424
r165 98 123 0.551426
r166 98 99 4.58464
r167 96 131 1.16709
r168 94 123 0.551426
r169 94 96 7.25207
r170 93 122 0.326018
r171 92 124 0.494161
r172 92 93 10.1279
r173 88 120 0.0828784
r174 88 90 1.82344
r175 86 125 0.494161
r176 86 87 15.8795
r177 85 122 0.326018
r178 84 120 0.551426
r179 84 85 15.5878
r180 83 120 0.551426
r181 82 87 0.652036
r182 82 83 4.58464
r183 74 118 1.16709
r184 69 102 1.16709
r185 65 90 1.16709
r186 56 145 0.0476429
r187 54 56 1.45875
r188 53 57 0.652036
r189 53 56 1.45875
r190 49 54 0.652036
r191 44 140 0.0476429
r192 42 44 1.45875
r193 41 45 0.652036
r194 41 44 1.45875
r195 37 42 0.652036
r196 32 131 0.238214
r197 30 32 1.45875
r198 29 33 0.652036
r199 29 32 1.45875
r200 25 30 0.652036
r201 11 57 3.8511
r202 11 49 3.8511
r203 10 74 0.185659
r204 8 69 0.185659
r205 5 45 3.8511
r206 5 37 3.8511
r207 3 33 3.1509
r208 3 25 3.1509
r209 2 65 0.185659
.ends

.subckt PM_G5_XNOR3_N2_C 2 4 6 8 20 23 32 40 43 47 52 57 67 86 94 100 Vss
c51 100 Vss 3.07518e-19
c52 94 Vss 0.00534351f
c53 86 Vss 0.010496f
c54 67 Vss 0.00399096f
c55 57 Vss 0.00459151f
c56 52 Vss 0.00198824f
c57 47 Vss 0.00148308f
c58 43 Vss 0.00113252f
c59 32 Vss 0.00492048f
c60 23 Vss 9.8832e-20
c61 20 Vss 0.221837f
c62 17 Vss 0.126125f
c63 15 Vss 0.0247918f
c64 4 Vss 0.133869f
r65 95 100 0.494161
r66 94 96 0.652036
r67 94 95 10.3363
r68 90 100 0.128424
r69 86 100 0.494161
r70 57 60 0.05
r71 52 67 1.16709
r72 52 96 2.37568
r73 47 90 2.45904
r74 43 60 1.16709
r75 43 86 25.2989
r76 40 43 0.0364688
r77 37 67 0.1
r78 32 47 1.16709
r79 23 57 0.0476429
r80 21 23 0.326018
r81 21 23 0.1167
r82 20 24 0.652036
r83 20 23 6.7686
r84 17 57 0.357321
r85 15 23 0.326018
r86 15 17 0.40845
r87 8 37 0.185659
r88 6 32 0.185659
r89 4 24 3.8511
r90 2 17 3.44265
.ends

.subckt PM_G5_XNOR3_N2_VSS 1 4 6 7 9 12 29 32 41 42 53 54 56 66 70 79 84 89 94
+ 99 102 105 114 119 128 130 131 132 137 138 143 151 159 160 161 Vss
c126 161 Vss 3.75522e-19
c127 160 Vss 3.88979e-19
c128 159 Vss 4.4306e-19
c129 143 Vss 0.00346584f
c130 138 Vss 8.41415e-19
c131 137 Vss 0.00629302f
c132 132 Vss 8.38477e-19
c133 131 Vss 0.00556756f
c134 130 Vss 0.00421531f
c135 128 Vss 0.00274186f
c136 119 Vss 0.00392167f
c137 114 Vss 0.00408379f
c138 105 Vss 0.00489622f
c139 102 Vss 0.00348146f
c140 99 Vss 0.00311148f
c141 94 Vss 7.25701e-19
c142 89 Vss 9.96742e-19
c143 84 Vss 0.00258358f
c144 79 Vss 0.00309974f
c145 70 Vss 0.00527641f
c146 66 Vss 0.00738563f
c147 56 Vss 1.02723e-19
c148 54 Vss 0.0347733f
c149 53 Vss 0.0999357f
c150 42 Vss 0.035088f
c151 41 Vss 0.0994129f
c152 32 Vss 9.8832e-20
c153 30 Vss 0.0348822f
c154 29 Vss 0.10032f
c155 9 Vss 0.270154f
c156 7 Vss 0.269158f
c157 6 Vss 0.00143442f
c158 1 Vss 0.232685f
r159 149 161 0.494161
r160 149 151 6.54354
r161 145 161 0.128424
r162 144 160 0.494161
r163 143 155 0.652036
r164 143 144 7.46046
r165 139 160 0.128424
r166 137 161 0.494161
r167 137 138 15.8795
r168 133 159 0.0828784
r169 131 160 0.494161
r170 131 132 13.0037
r171 130 138 0.652036
r172 129 159 0.551426
r173 129 130 12.5036
r174 128 159 0.551426
r175 127 132 0.652036
r176 127 128 7.66886
r177 102 151 1.50043
r178 99 102 5.835
r179 94 119 1.16709
r180 94 155 2.16729
r181 89 114 1.16709
r182 89 145 2.16729
r183 84 139 5.2515
r184 79 105 1.16709
r185 79 133 4.33978
r186 70 99 1.16709
r187 66 84 1.16709
r188 56 119 0.0476429
r189 54 56 1.45875
r190 53 57 0.652036
r191 53 56 1.45875
r192 49 54 0.652036
r193 44 114 0.0476429
r194 42 44 1.45875
r195 41 45 0.652036
r196 41 44 1.45875
r197 37 42 0.652036
r198 32 105 0.238214
r199 30 32 1.45875
r200 29 33 0.652036
r201 29 32 1.45875
r202 25 30 0.652036
r203 12 70 0.185659
r204 9 57 3.8511
r205 9 49 3.8511
r206 7 45 3.8511
r207 7 37 3.8511
r208 6 66 0.185659
r209 4 66 0.185659
r210 1 33 3.1509
r211 1 25 3.1509
.ends

.subckt PM_G5_XNOR3_N2_CI 2 4 6 8 23 26 31 34 39 44 79 80 85 91 Vss
c48 91 Vss 2.53341e-19
c49 85 Vss 0.00608182f
c50 80 Vss 3.61784e-19
c51 79 Vss 0.00606729f
c52 44 Vss 0.00187346f
c53 39 Vss 0.00150573f
c54 34 Vss 0.00581447f
c55 31 Vss 0.00501461f
c56 26 Vss 0.00386883f
c57 23 Vss 0.00546807f
c58 4 Vss 0.00143442f
r59 86 91 0.441572
r60 85 87 0.655813
r61 85 86 9.04425
r62 81 91 0.174814
r63 79 91 0.441572
r64 79 80 19.1096
r65 75 80 0.655813
r66 44 87 2.41736
r67 39 81 2.41736
r68 34 75 13.4205
r69 31 44 1.16709
r70 26 39 1.16709
r71 23 34 1.16709
r72 8 31 0.185659
r73 6 26 0.185659
r74 4 23 0.185659
r75 2 23 0.185659
.ends

.subckt PM_G5_XNOR3_N2_A 2 4 5 7 20 44 45 49 55 58 60 61 66 69 70 73 78 Vss
c79 78 Vss 0.00548899f
c80 73 Vss 0.00489228f
c81 70 Vss 0.00566456f
c82 69 Vss 4.97253e-19
c83 61 Vss 5.64597e-19
c84 60 Vss 6.06847e-19
c85 58 Vss 0.00443885f
c86 55 Vss 0.00696223f
c87 49 Vss 0.135055f
c88 45 Vss 0.127825f
c89 44 Vss 9.8832e-20
c90 20 Vss 0.21515f
c91 17 Vss 0.129208f
c92 15 Vss 0.0247918f
c93 5 Vss 1.22081f
c94 4 Vss 0.139574f
r95 78 81 0.05
r96 69 81 1.16709
r97 69 70 0.531835
r98 64 73 1.16709
r99 64 66 0.125036
r100 61 64 0.833571
r101 60 70 10.4613
r102 57 60 0.652036
r103 57 58 8.66914
r104 56 61 0.0685365
r105 55 58 0.652036
r106 55 56 10.2113
r107 47 49 4.53833
r108 44 78 0.0238214
r109 44 45 2.26917
r110 41 44 2.26917
r111 34 49 0.00605528
r112 33 45 0.00605528
r113 28 47 0.00605528
r114 27 41 0.00605528
r115 23 73 0.0952857
r116 21 23 0.326018
r117 21 23 0.1167
r118 20 24 0.652036
r119 20 23 6.7686
r120 17 23 0.3335
r121 15 23 0.326018
r122 15 17 0.2334
r123 7 34 3.8511
r124 7 28 3.8511
r125 5 7 15.4044
r126 5 33 3.8511
r127 5 7 15.4044
r128 5 27 3.8511
r129 4 24 3.8511
r130 2 17 3.6177
.ends

.subckt PM_G5_XNOR3_N2_BI 2 4 6 8 16 23 29 32 37 42 51 56 64 65 71 77 82 83 Vss
c69 83 Vss 1.50773e-19
c70 82 Vss 0.00211439f
c71 77 Vss 0.00104035f
c72 71 Vss 3.29809e-19
c73 65 Vss 2.46443e-19
c74 64 Vss 0.00335376f
c75 56 Vss 0.00250661f
c76 51 Vss 0.00216609f
c77 42 Vss 0.00132272f
c78 37 Vss 9.45807e-19
c79 32 Vss 0.00229686f
c80 29 Vss 0.00450667f
c81 23 Vss 1.05854e-19
c82 16 Vss 0.111942f
c83 8 Vss 0.111942f
c84 4 Vss 0.00143442f
r85 81 83 0.65409
r86 81 82 3.42052
r87 77 82 0.652979
r88 64 71 0.0685365
r89 64 65 13.2121
r90 60 65 0.652036
r91 42 56 1.16709
r92 42 83 2.00578
r93 37 51 1.16709
r94 37 77 2.03284
r95 37 71 2.08393
r96 32 60 5.2515
r97 29 32 1.16709
r98 23 56 0.50025
r99 16 51 0.50025
r100 8 23 3.09255
r101 6 16 3.09255
r102 4 29 0.185659
r103 2 29 0.185659
.ends

.subckt PM_G5_XNOR3_N2_AI 2 4 5 7 31 37 43 50 55 64 72 Vss
c47 72 Vss 2.58509e-19
c48 64 Vss 0.005486f
c49 55 Vss 0.0041561f
c50 50 Vss 8.67602e-19
c51 43 Vss 0.00448756f
c52 37 Vss 0.127877f
c53 31 Vss 0.131783f
c54 5 Vss 1.2083f
c55 4 Vss 0.00143442f
r56 68 72 0.655813
r57 55 64 1.16709
r58 55 72 12.0347
r59 50 68 2.41736
r60 43 50 1.16709
r61 36 64 0.0238214
r62 36 37 2.334
r63 33 36 2.20433
r64 29 31 4.53833
r65 24 37 0.00605528
r66 23 31 0.00605528
r67 18 33 0.00605528
r68 17 29 0.00605528
r69 7 24 3.8511
r70 7 18 3.8511
r71 5 7 15.4044
r72 5 23 3.8511
r73 5 7 15.4044
r74 5 17 3.8511
r75 4 43 0.185659
r76 2 43 0.185659
.ends

.subckt PM_G5_XNOR3_N2_B 2 4 6 8 16 17 24 28 31 42 45 50 55 60 65 69 74 75 82
+ Vss
c65 82 Vss 3.53127e-19
c66 75 Vss 3.16204e-19
c67 74 Vss 7.66068e-19
c68 69 Vss 0.00368257f
c69 65 Vss 0.00255458f
c70 60 Vss 0.0023582f
c71 55 Vss 0.00157585f
c72 50 Vss 0.00115924f
c73 45 Vss 7.04295e-20
c74 42 Vss 5.36415e-19
c75 31 Vss 0.111942f
c76 24 Vss 1.02723e-19
c77 20 Vss 0.0247918f
c78 17 Vss 0.0338452f
c79 16 Vss 0.183686f
c80 6 Vss 0.112114f
c81 4 Vss 0.122719f
c82 2 Vss 0.13381f
r83 74 75 0.65409
r84 73 74 3.38028
r85 69 73 0.65409
r86 50 65 1.16709
r87 50 75 2.00578
r88 45 60 1.16709
r89 45 69 1.96931
r90 45 82 9.55481
r91 38 55 1.16709
r92 38 82 0.4602
r93 38 42 0.145875
r94 36 55 0.309679
r95 31 65 0.50025
r96 28 60 0.50025
r97 24 55 0.214393
r98 20 36 0.326018
r99 20 24 0.75855
r100 17 36 6.7686
r101 16 36 0.326018
r102 16 36 0.1167
r103 13 17 0.652036
r104 8 31 3.09255
r105 6 28 3.09255
r106 4 24 3.09255
r107 2 13 3.8511
.ends

.subckt PM_G5_XNOR3_N2_Z 2 4 6 8 23 27 30 33 Vss
c29 30 Vss 0.00359454f
c30 27 Vss 0.00857889f
c31 23 Vss 0.0074536f
c32 8 Vss 0.00143442f
c33 6 Vss 0.00143442f
r34 33 35 5.50157
r35 30 33 5.50157
r36 27 35 1.16709
r37 23 30 1.16709
r38 8 27 0.185659
r39 6 23 0.185659
r40 4 27 0.185659
r41 2 23 0.185659
.ends

.subckt G5_XNOR3_N2  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI13.X0 N_CI_XI13.X0_D N_VSS_XI13.X0_PGD N_C_XI13.X0_CG N_VSS_XI13.X0_PGD
+ N_VDD_XI13.X0_S TIGFET_HPNW8
XI16.X0 N_CI_XI16.X0_D N_VDD_XI16.X0_PGD N_C_XI16.X0_CG N_VDD_XI16.X0_PGD
+ N_VSS_XI16.X0_S TIGFET_HPNW8
XI15.X0 N_BI_XI15.X0_D N_VDD_XI15.X0_PGD N_B_XI15.X0_CG N_VDD_XI15.X0_PGD
+ N_VSS_XI15.X0_S TIGFET_HPNW8
XI11.X0 N_AI_XI11.X0_D N_VSS_XI11.X0_PGD N_A_XI11.X0_CG N_VSS_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW8
XI12.X0 N_BI_XI12.X0_D N_VSS_XI12.X0_PGD N_B_XI12.X0_CG N_VSS_XI12.X0_PGD
+ N_VDD_XI12.X0_S TIGFET_HPNW8
XI14.X0 N_AI_XI14.X0_D N_VDD_XI14.X0_PGD N_A_XI14.X0_CG N_VDD_XI14.X0_PGD
+ N_VSS_XI14.X0_S TIGFET_HPNW8
XI19.X0 N_Z_XI19.X0_D N_AI_XI19.X0_PGD N_B_XI19.X0_CG N_AI_XI19.X0_PGD
+ N_C_XI19.X0_S TIGFET_HPNW8
XI17.X0 N_Z_XI17.X0_D N_AI_XI17.X0_PGD N_BI_XI17.X0_CG N_AI_XI17.X0_PGD
+ N_CI_XI17.X0_S TIGFET_HPNW8
XI20.X0 N_Z_XI20.X0_D N_A_XI20.X0_PGD N_BI_XI20.X0_CG N_A_XI20.X0_PGD
+ N_C_XI20.X0_S TIGFET_HPNW8
XI18.X0 N_Z_XI18.X0_D N_A_XI18.X0_PGD N_B_XI18.X0_CG N_A_XI18.X0_PGD
+ N_CI_XI18.X0_S TIGFET_HPNW8
*
x_PM_G5_XNOR3_N2_VDD N_VDD_XI13.X0_S N_VDD_XI16.X0_PGD N_VDD_XI15.X0_PGD
+ N_VDD_XI11.X0_S N_VDD_XI12.X0_S N_VDD_XI14.X0_PGD N_VDD_c_115_p N_VDD_c_20_p
+ N_VDD_c_25_p N_VDD_c_3_p N_VDD_c_95_p N_VDD_c_106_p N_VDD_c_21_p N_VDD_c_77_p
+ N_VDD_c_107_p N_VDD_c_5_p N_VDD_c_6_p N_VDD_c_13_p N_VDD_c_4_p N_VDD_c_65_p
+ N_VDD_c_30_p N_VDD_c_66_p N_VDD_c_31_p N_VDD_c_17_p N_VDD_c_67_p N_VDD_c_22_p
+ N_VDD_c_10_p N_VDD_c_26_p N_VDD_c_38_p N_VDD_c_11_p N_VDD_c_61_p VDD
+ N_VDD_c_69_p N_VDD_c_73_p N_VDD_c_32_p N_VDD_c_43_p N_VDD_c_39_p Vss
+ PM_G5_XNOR3_N2_VDD
x_PM_G5_XNOR3_N2_C N_C_XI13.X0_CG N_C_XI16.X0_CG N_C_XI19.X0_S N_C_XI20.X0_S
+ N_C_c_118_n N_C_c_129_p N_C_c_121_n C N_C_c_122_n N_C_c_147_p N_C_c_144_p
+ N_C_c_124_n N_C_c_165_p N_C_c_126_n N_C_c_149_p N_C_c_154_p Vss
+ PM_G5_XNOR3_N2_C
x_PM_G5_XNOR3_N2_VSS N_VSS_XI13.X0_PGD N_VSS_XI16.X0_S N_VSS_XI15.X0_S
+ N_VSS_XI11.X0_PGD N_VSS_XI12.X0_PGD N_VSS_XI14.X0_S N_VSS_c_176_n
+ N_VSS_c_234_n N_VSS_c_177_n N_VSS_c_179_n N_VSS_c_180_n N_VSS_c_181_n
+ N_VSS_c_288_p N_VSS_c_183_n N_VSS_c_249_p N_VSS_c_184_n N_VSS_c_189_n
+ N_VSS_c_192_n N_VSS_c_196_n N_VSS_c_200_n N_VSS_c_203_n N_VSS_c_204_n
+ N_VSS_c_207_n N_VSS_c_211_n N_VSS_c_215_n N_VSS_c_218_n N_VSS_c_220_n
+ N_VSS_c_221_n N_VSS_c_222_n N_VSS_c_226_n N_VSS_c_227_n VSS N_VSS_c_230_n
+ N_VSS_c_231_n N_VSS_c_232_n Vss PM_G5_XNOR3_N2_VSS
x_PM_G5_XNOR3_N2_CI N_CI_XI13.X0_D N_CI_XI16.X0_D N_CI_XI17.X0_S N_CI_XI18.X0_S
+ N_CI_c_294_n N_CI_c_306_n N_CI_c_336_p N_CI_c_295_n N_CI_c_314_n N_CI_c_303_n
+ N_CI_c_299_n N_CI_c_319_n N_CI_c_322_p N_CI_c_331_p Vss PM_G5_XNOR3_N2_CI
x_PM_G5_XNOR3_N2_A N_A_XI11.X0_CG N_A_XI14.X0_CG N_A_XI20.X0_PGD N_A_XI18.X0_PGD
+ N_A_c_342_n N_A_c_376_p N_A_c_392_p N_A_c_394_p N_A_c_343_n N_A_c_349_n
+ N_A_c_350_n N_A_c_351_n A N_A_c_360_n N_A_c_361_n N_A_c_353_n N_A_c_382_p Vss
+ PM_G5_XNOR3_N2_A
x_PM_G5_XNOR3_N2_BI N_BI_XI15.X0_D N_BI_XI12.X0_D N_BI_XI17.X0_CG
+ N_BI_XI20.X0_CG N_BI_c_456_p N_BI_c_443_n N_BI_c_421_n N_BI_c_423_n
+ N_BI_c_459_p N_BI_c_438_n N_BI_c_457_p N_BI_c_450_n N_BI_c_427_n N_BI_c_454_n
+ N_BI_c_455_n N_BI_c_430_n N_BI_c_482_p N_BI_c_431_n Vss PM_G5_XNOR3_N2_BI
x_PM_G5_XNOR3_N2_AI N_AI_XI11.X0_D N_AI_XI14.X0_D N_AI_XI19.X0_PGD
+ N_AI_XI17.X0_PGD N_AI_c_499_n N_AI_c_491_n N_AI_c_492_n N_AI_c_494_n
+ N_AI_c_497_n N_AI_c_506_n N_AI_c_507_n Vss PM_G5_XNOR3_N2_AI
x_PM_G5_XNOR3_N2_B N_B_XI15.X0_CG N_B_XI12.X0_CG N_B_XI19.X0_CG N_B_XI18.X0_CG
+ N_B_c_538_n N_B_c_539_n N_B_c_545_n N_B_c_558_n N_B_c_559_n B N_B_c_562_n
+ N_B_c_551_n N_B_c_548_n N_B_c_567_n N_B_c_568_n N_B_c_540_n N_B_c_588_n
+ N_B_c_552_n N_B_c_550_n Vss PM_G5_XNOR3_N2_B
x_PM_G5_XNOR3_N2_Z N_Z_XI19.X0_D N_Z_XI17.X0_D N_Z_XI20.X0_D N_Z_XI18.X0_D
+ N_Z_c_602_n N_Z_c_608_n N_Z_c_606_n Z Vss PM_G5_XNOR3_N2_Z
cc_1 N_VDD_XI15.X0_PGD N_C_XI16.X0_CG 0.00111638f
cc_2 N_VDD_XI16.X0_PGD N_C_c_118_n 4.18107e-19
cc_3 N_VDD_c_3_p N_C_c_118_n 0.00111638f
cc_4 N_VDD_c_4_p N_C_c_118_n 0.00134502f
cc_5 N_VDD_c_5_p N_C_c_121_n 3.43419e-19
cc_6 N_VDD_c_6_p N_C_c_122_n 4.34606e-19
cc_7 N_VDD_c_4_p N_C_c_122_n 0.00156986f
cc_8 N_VDD_c_6_p N_C_c_124_n 4.60895e-19
cc_9 N_VDD_c_4_p N_C_c_124_n 2.85335e-19
cc_10 N_VDD_c_10_p N_C_c_126_n 4.68396e-19
cc_11 N_VDD_c_11_p N_C_c_126_n 7.76004e-19
cc_12 N_VDD_XI16.X0_PGD N_VSS_XI13.X0_PGD 0.00162006f
cc_13 N_VDD_c_13_p N_VSS_XI13.X0_PGD 2.10457e-19
cc_14 N_VDD_c_4_p N_VSS_XI13.X0_PGD 2.00345e-19
cc_15 N_VDD_XI15.X0_PGD N_VSS_XI11.X0_PGD 2.37403e-19
cc_16 N_VDD_XI14.X0_PGD N_VSS_XI11.X0_PGD 0.00200476f
cc_17 N_VDD_c_17_p N_VSS_XI11.X0_PGD 2.94729e-19
cc_18 N_VDD_XI15.X0_PGD N_VSS_XI12.X0_PGD 0.00200584f
cc_19 N_VDD_XI14.X0_PGD N_VSS_XI12.X0_PGD 2.24644e-19
cc_20 N_VDD_c_20_p N_VSS_c_176_n 0.00162006f
cc_21 N_VDD_c_21_p N_VSS_c_177_n 0.00200476f
cc_22 N_VDD_c_22_p N_VSS_c_177_n 2.84318e-19
cc_23 N_VDD_c_22_p N_VSS_c_179_n 3.9313e-19
cc_24 N_VDD_c_11_p N_VSS_c_180_n 2.35523e-19
cc_25 N_VDD_c_25_p N_VSS_c_181_n 0.00200584f
cc_26 N_VDD_c_26_p N_VSS_c_181_n 3.9313e-19
cc_27 N_VDD_c_4_p N_VSS_c_183_n 3.4118e-19
cc_28 N_VDD_c_13_p N_VSS_c_184_n 4.32468e-19
cc_29 N_VDD_c_4_p N_VSS_c_184_n 4.11891e-19
cc_30 N_VDD_c_30_p N_VSS_c_184_n 0.00126261f
cc_31 N_VDD_c_31_p N_VSS_c_184_n 3.98949e-19
cc_32 N_VDD_c_32_p N_VSS_c_184_n 3.48267e-19
cc_33 N_VDD_c_4_p N_VSS_c_189_n 3.98099e-19
cc_34 N_VDD_c_10_p N_VSS_c_189_n 7.41581e-19
cc_35 N_VDD_c_11_p N_VSS_c_189_n 5.12345e-19
cc_36 N_VDD_c_17_p N_VSS_c_192_n 6.9475e-19
cc_37 N_VDD_c_22_p N_VSS_c_192_n 0.00161703f
cc_38 N_VDD_c_38_p N_VSS_c_192_n 9.10421e-19
cc_39 N_VDD_c_39_p N_VSS_c_192_n 3.48267e-19
cc_40 N_VDD_c_10_p N_VSS_c_196_n 6.80981e-19
cc_41 N_VDD_c_26_p N_VSS_c_196_n 0.00161703f
cc_42 N_VDD_c_11_p N_VSS_c_196_n 0.00260511f
cc_43 N_VDD_c_43_p N_VSS_c_196_n 3.48267e-19
cc_44 N_VDD_XI14.X0_PGD N_VSS_c_200_n 2.99706e-19
cc_45 N_VDD_c_38_p N_VSS_c_200_n 0.00524008f
cc_46 N_VDD_c_39_p N_VSS_c_200_n 9.58524e-19
cc_47 N_VDD_c_22_p N_VSS_c_203_n 0.00398219f
cc_48 N_VDD_c_13_p N_VSS_c_204_n 4.41003e-19
cc_49 N_VDD_c_31_p N_VSS_c_204_n 3.89161e-19
cc_50 N_VDD_c_32_p N_VSS_c_204_n 6.39485e-19
cc_51 N_VDD_c_17_p N_VSS_c_207_n 3.48267e-19
cc_52 N_VDD_c_22_p N_VSS_c_207_n 2.26455e-19
cc_53 N_VDD_c_38_p N_VSS_c_207_n 3.99794e-19
cc_54 N_VDD_c_39_p N_VSS_c_207_n 6.489e-19
cc_55 N_VDD_c_10_p N_VSS_c_211_n 3.82294e-19
cc_56 N_VDD_c_26_p N_VSS_c_211_n 2.26455e-19
cc_57 N_VDD_c_11_p N_VSS_c_211_n 9.55109e-19
cc_58 N_VDD_c_43_p N_VSS_c_211_n 6.46219e-19
cc_59 N_VDD_c_6_p N_VSS_c_215_n 0.00346699f
cc_60 N_VDD_c_13_p N_VSS_c_215_n 0.0014056f
cc_61 N_VDD_c_61_p N_VSS_c_215_n 0.0010705f
cc_62 N_VDD_c_13_p N_VSS_c_218_n 0.00935412f
cc_63 N_VDD_c_31_p N_VSS_c_218_n 0.00107899f
cc_64 N_VDD_c_4_p N_VSS_c_220_n 0.00942626f
cc_65 N_VDD_c_65_p N_VSS_c_221_n 0.00107364f
cc_66 N_VDD_c_66_p N_VSS_c_222_n 0.00824191f
cc_67 N_VDD_c_67_p N_VSS_c_222_n 7.27535e-19
cc_68 N_VDD_c_22_p N_VSS_c_222_n 0.00364308f
cc_69 N_VDD_c_69_p N_VSS_c_222_n 0.00146091f
cc_70 N_VDD_c_13_p N_VSS_c_226_n 0.00107577f
cc_71 N_VDD_c_4_p N_VSS_c_227_n 0.00143205f
cc_72 N_VDD_c_26_p N_VSS_c_227_n 0.00595362f
cc_73 N_VDD_c_73_p N_VSS_c_227_n 0.00107225f
cc_74 N_VDD_c_13_p N_VSS_c_230_n 0.00112682f
cc_75 N_VDD_c_4_p N_VSS_c_231_n 0.00107375f
cc_76 N_VDD_c_22_p N_VSS_c_232_n 7.74609e-19
cc_77 N_VDD_c_77_p N_CI_c_294_n 3.43419e-19
cc_78 N_VDD_c_77_p N_CI_c_295_n 3.48267e-19
cc_79 N_VDD_c_4_p N_CI_c_295_n 4.34701e-19
cc_80 N_VDD_c_30_p N_CI_c_295_n 5.61123e-19
cc_81 N_VDD_c_31_p N_CI_c_295_n 0.00251349f
cc_82 N_VDD_c_17_p N_CI_c_299_n 9.69348e-19
cc_83 N_VDD_c_67_p N_CI_c_299_n 5.49852e-19
cc_84 N_VDD_XI14.X0_PGD N_A_c_342_n 3.94724e-19
cc_85 N_VDD_XI14.X0_PGD N_A_c_343_n 4.9801e-19
cc_86 N_VDD_c_5_p N_A_c_343_n 2.69869e-19
cc_87 N_VDD_c_22_p N_A_c_343_n 2.92916e-19
cc_88 N_VDD_c_38_p N_A_c_343_n 2.57998e-19
cc_89 N_VDD_c_11_p N_A_c_343_n 3.18391e-19
cc_90 N_VDD_c_39_p N_A_c_343_n 4.99558e-19
cc_91 N_VDD_c_5_p N_A_c_349_n 9.18655e-19
cc_92 N_VDD_c_11_p N_A_c_350_n 0.00561464f
cc_93 N_VDD_c_31_p N_A_c_351_n 0.00109781f
cc_94 N_VDD_c_10_p N_A_c_351_n 2.35756e-19
cc_95 N_VDD_c_95_p N_A_c_353_n 3.65048e-19
cc_96 N_VDD_c_31_p N_A_c_353_n 5.7233e-19
cc_97 N_VDD_c_43_p N_A_c_353_n 2.01103e-19
cc_98 N_VDD_c_5_p N_BI_c_421_n 3.43419e-19
cc_99 N_VDD_c_11_p N_BI_c_421_n 3.48267e-19
cc_100 N_VDD_c_5_p N_BI_c_423_n 3.48267e-19
cc_101 N_VDD_c_31_p N_BI_c_423_n 9.37844e-19
cc_102 N_VDD_c_26_p N_BI_c_423_n 4.34701e-19
cc_103 N_VDD_c_11_p N_BI_c_423_n 4.99861e-19
cc_104 N_VDD_c_26_p N_BI_c_427_n 2.93466e-19
cc_105 N_VDD_XI14.X0_PGD N_AI_XI19.X0_PGD 3.10667e-19
cc_106 N_VDD_c_106_p N_AI_c_491_n 3.10667e-19
cc_107 N_VDD_c_107_p N_AI_c_492_n 3.43419e-19
cc_108 N_VDD_c_67_p N_AI_c_492_n 3.73302e-19
cc_109 N_VDD_c_107_p N_AI_c_494_n 3.48267e-19
cc_110 N_VDD_c_67_p N_AI_c_494_n 5.23123e-19
cc_111 N_VDD_c_22_p N_AI_c_494_n 4.34701e-19
cc_112 N_VDD_c_38_p N_AI_c_497_n 0.00114561f
cc_113 N_VDD_XI16.X0_PGD N_B_XI15.X0_CG 8.43351e-19
cc_114 N_VDD_XI15.X0_PGD N_B_c_538_n 3.99339e-19
cc_115 N_VDD_c_115_p N_B_c_539_n 8.43351e-19
cc_116 N_VDD_c_11_p N_B_c_540_n 4.93279e-19
cc_117 N_C_c_118_n N_VSS_XI13.X0_PGD 4.18107e-19
cc_118 N_C_c_129_p N_VSS_c_234_n 9.69352e-19
cc_119 N_C_c_122_n N_VSS_c_184_n 7.02166e-19
cc_120 N_C_c_124_n N_VSS_c_184_n 3.26762e-19
cc_121 N_C_c_122_n N_VSS_c_189_n 2.08725e-19
cc_122 N_C_c_126_n N_VSS_c_189_n 0.00161414f
cc_123 N_C_c_126_n N_VSS_c_196_n 0.00142183f
cc_124 N_C_c_122_n N_VSS_c_204_n 3.26762e-19
cc_125 N_C_c_124_n N_VSS_c_204_n 2.75266e-19
cc_126 N_C_c_122_n N_VSS_c_215_n 4.20305e-19
cc_127 N_C_c_126_n N_VSS_c_215_n 2.33946e-19
cc_128 N_C_c_122_n N_VSS_c_220_n 0.00170504f
cc_129 N_C_c_126_n N_VSS_c_220_n 0.00306503f
cc_130 N_C_c_126_n N_VSS_c_227_n 0.00185247f
cc_131 N_C_c_118_n N_CI_c_294_n 6.55689e-19
cc_132 N_C_c_126_n N_CI_c_295_n 0.00101197f
cc_133 N_C_c_144_p N_CI_c_303_n 2.42706e-19
cc_134 N_C_c_126_n N_A_c_343_n 3.07864e-19
cc_135 N_C_c_121_n N_A_c_349_n 8.20481e-19
cc_136 N_C_c_147_p N_A_c_349_n 0.00174813f
cc_137 N_C_c_126_n N_A_c_350_n 3.74205e-19
cc_138 N_C_c_149_p N_A_c_360_n 3.98753e-19
cc_139 N_C_c_121_n N_A_c_361_n 8.20481e-19
cc_140 N_C_c_147_p N_A_c_361_n 0.00170439f
cc_141 N_C_c_126_n N_A_c_361_n 3.354e-19
cc_142 N_C_c_149_p N_A_c_361_n 0.00192636f
cc_143 N_C_c_154_p N_A_c_361_n 2.01694e-19
cc_144 N_C_c_126_n N_BI_c_423_n 4.79207e-19
cc_145 N_C_c_126_n N_BI_c_427_n 5.14704e-19
cc_146 N_C_c_149_p N_BI_c_430_n 5.49277e-19
cc_147 N_C_c_149_p N_BI_c_431_n 0.00181681f
cc_148 N_C_c_147_p N_B_c_540_n 0.00168209f
cc_149 N_C_c_126_n N_B_c_540_n 0.00270379f
cc_150 N_C_c_149_p N_B_c_540_n 0.0010597f
cc_151 N_C_c_121_n N_Z_c_602_n 3.43419e-19
cc_152 N_C_c_147_p N_Z_c_602_n 3.48267e-19
cc_153 N_C_c_144_p N_Z_c_602_n 3.48267e-19
cc_154 N_C_c_165_p N_Z_c_602_n 3.43419e-19
cc_155 N_C_c_147_p N_Z_c_606_n 6.10113e-19
cc_156 N_C_c_144_p N_Z_c_606_n 5.74072e-19
cc_157 N_VSS_c_183_n N_CI_c_294_n 3.43419e-19
cc_158 N_VSS_c_189_n N_CI_c_294_n 3.48267e-19
cc_159 N_VSS_c_249_p N_CI_c_306_n 3.43419e-19
cc_160 N_VSS_c_200_n N_CI_c_306_n 3.48267e-19
cc_161 N_VSS_c_183_n N_CI_c_295_n 3.48267e-19
cc_162 N_VSS_c_184_n N_CI_c_295_n 5.78167e-19
cc_163 N_VSS_c_189_n N_CI_c_295_n 0.00107566f
cc_164 N_VSS_c_215_n N_CI_c_295_n 3.18991e-19
cc_165 N_VSS_c_218_n N_CI_c_295_n 0.00247956f
cc_166 N_VSS_c_220_n N_CI_c_295_n 2.82247e-19
cc_167 N_VSS_c_249_p N_CI_c_314_n 3.48267e-19
cc_168 N_VSS_c_200_n N_CI_c_314_n 9.64594e-19
cc_169 N_VSS_c_192_n N_CI_c_299_n 0.00118348f
cc_170 N_VSS_c_203_n N_CI_c_299_n 0.0033401f
cc_171 N_VSS_c_222_n N_CI_c_299_n 2.16087e-19
cc_172 N_VSS_c_222_n N_CI_c_319_n 0.00291606f
cc_173 N_VSS_XI11.X0_PGD N_A_c_342_n 3.91527e-19
cc_174 N_VSS_c_249_p N_A_c_343_n 5.38503e-19
cc_175 N_VSS_c_200_n N_A_c_343_n 8.92829e-19
cc_176 N_VSS_c_203_n N_A_c_343_n 2.86582e-19
cc_177 N_VSS_c_192_n N_A_c_351_n 3.11664e-19
cc_178 N_VSS_c_207_n N_A_c_351_n 3.1261e-19
cc_179 N_VSS_c_192_n N_A_c_353_n 3.04912e-19
cc_180 N_VSS_c_207_n N_A_c_353_n 0.00110478f
cc_181 N_VSS_c_183_n N_BI_c_421_n 3.43419e-19
cc_182 N_VSS_c_189_n N_BI_c_421_n 3.48267e-19
cc_183 N_VSS_c_183_n N_BI_c_423_n 3.48267e-19
cc_184 N_VSS_c_189_n N_BI_c_423_n 0.00102079f
cc_185 N_VSS_c_227_n N_BI_c_423_n 2.89128e-19
cc_186 N_VSS_XI12.X0_PGD N_AI_XI19.X0_PGD 2.79882e-19
cc_187 N_VSS_c_180_n N_AI_c_499_n 2.79882e-19
cc_188 N_VSS_c_249_p N_AI_c_492_n 3.43419e-19
cc_189 N_VSS_c_200_n N_AI_c_492_n 3.48267e-19
cc_190 N_VSS_c_249_p N_AI_c_494_n 3.48267e-19
cc_191 N_VSS_c_200_n N_AI_c_494_n 0.001398f
cc_192 N_VSS_c_200_n N_AI_c_497_n 0.00172519f
cc_193 N_VSS_c_203_n N_AI_c_497_n 0.00643151f
cc_194 N_VSS_c_200_n N_AI_c_506_n 2.82216e-19
cc_195 N_VSS_c_192_n N_AI_c_507_n 0.00195338f
cc_196 N_VSS_c_203_n N_AI_c_507_n 0.00167155f
cc_197 N_VSS_XI12.X0_PGD N_B_c_538_n 3.96142e-19
cc_198 N_VSS_c_288_p N_B_c_545_n 0.00112923f
cc_199 N_VSS_c_196_n B 3.70276e-19
cc_200 N_VSS_c_211_n B 3.65807e-19
cc_201 N_VSS_c_196_n N_B_c_548_n 3.65807e-19
cc_202 N_VSS_c_211_n N_B_c_548_n 3.61194e-19
cc_203 N_VSS_c_196_n N_B_c_550_n 4.74612e-19
cc_204 N_CI_c_299_n N_A_c_343_n 4.46962e-19
cc_205 N_CI_c_295_n N_BI_c_423_n 0.00125164f
cc_206 N_CI_c_322_p N_BI_c_438_n 6.43262e-19
cc_207 N_CI_c_314_n N_BI_c_427_n 5.16242e-19
cc_208 N_CI_c_299_n N_BI_c_427_n 0.00141805f
cc_209 N_CI_c_322_p N_BI_c_430_n 0.00184196f
cc_210 N_CI_c_295_n N_AI_c_494_n 5.9142e-19
cc_211 N_CI_c_314_n N_AI_c_494_n 5.87215e-19
cc_212 N_CI_c_314_n N_AI_c_497_n 0.00175375f
cc_213 N_CI_c_299_n N_AI_c_497_n 0.0058239f
cc_214 N_CI_c_322_p N_AI_c_497_n 0.00302067f
cc_215 N_CI_c_331_p N_AI_c_497_n 9.17939e-19
cc_216 N_CI_c_299_n N_AI_c_507_n 6.9086e-19
cc_217 N_CI_c_322_p N_B_c_551_n 8.97242e-19
cc_218 N_CI_c_322_p N_B_c_552_n 2.22052e-19
cc_219 N_CI_c_306_n N_Z_c_608_n 3.43419e-19
cc_220 N_CI_c_336_p N_Z_c_608_n 3.43419e-19
cc_221 N_CI_c_314_n N_Z_c_608_n 3.48267e-19
cc_222 N_CI_c_303_n N_Z_c_608_n 3.48267e-19
cc_223 N_CI_c_336_p N_Z_c_606_n 3.48267e-19
cc_224 N_CI_c_314_n N_Z_c_606_n 6.09821e-19
cc_225 N_CI_c_303_n N_Z_c_606_n 5.71987e-19
cc_226 N_A_XI20.X0_PGD N_BI_XI20.X0_CG 9.65637e-19
cc_227 N_A_c_376_p N_BI_c_443_n 9.50932e-19
cc_228 N_A_c_343_n N_BI_c_421_n 2.69869e-19
cc_229 N_A_c_343_n N_BI_c_423_n 2.84781e-19
cc_230 N_A_c_349_n N_BI_c_423_n 7.93978e-19
cc_231 N_A_c_360_n N_BI_c_438_n 5.59762e-19
cc_232 N_A_c_361_n N_BI_c_438_n 2.11253e-19
cc_233 N_A_c_382_p N_BI_c_438_n 3.26762e-19
cc_234 N_A_XI20.X0_PGD N_BI_c_450_n 0.00133285f
cc_235 N_A_c_382_p N_BI_c_450_n 2.75266e-19
cc_236 N_A_c_343_n N_BI_c_427_n 0.0032866f
cc_237 N_A_c_349_n N_BI_c_427_n 0.00143358f
cc_238 N_A_c_343_n N_BI_c_454_n 6.46327e-19
cc_239 N_A_c_343_n N_BI_c_455_n 2.29103e-19
cc_240 N_A_XI20.X0_PGD N_AI_XI19.X0_PGD 0.0174153f
cc_241 N_A_c_349_n N_AI_XI19.X0_PGD 9.9436e-19
cc_242 N_A_c_361_n N_AI_XI19.X0_PGD 0.00100436f
cc_243 N_A_c_392_p N_AI_c_499_n 0.00199603f
cc_244 N_A_c_361_n N_AI_c_499_n 0.001261f
cc_245 N_A_c_394_p N_AI_c_491_n 0.00201004f
cc_246 N_A_c_342_n N_AI_c_492_n 6.8653e-19
cc_247 N_A_c_343_n N_AI_c_494_n 8.04759e-19
cc_248 N_A_c_343_n N_AI_c_497_n 0.00144224f
cc_249 N_A_c_342_n N_B_c_538_n 0.00359928f
cc_250 N_A_c_343_n N_B_c_538_n 3.71868e-19
cc_251 N_A_c_351_n N_B_c_539_n 3.71868e-19
cc_252 N_A_c_353_n N_B_c_539_n 5.91713e-19
cc_253 N_A_c_343_n N_B_c_545_n 3.88197e-19
cc_254 N_A_c_361_n N_B_c_558_n 2.74063e-19
cc_255 N_A_XI20.X0_PGD N_B_c_559_n 9.65637e-19
cc_256 N_A_c_343_n B 7.21228e-19
cc_257 N_A_c_349_n B 4.92712e-19
cc_258 N_A_c_349_n N_B_c_562_n 3.80412e-19
cc_259 N_A_c_361_n N_B_c_562_n 3.68965e-19
cc_260 N_A_c_361_n N_B_c_551_n 4.34114e-19
cc_261 N_A_c_342_n N_B_c_548_n 6.98561e-19
cc_262 N_A_c_349_n N_B_c_548_n 6.04163e-19
cc_263 N_A_c_349_n N_B_c_567_n 3.37713e-19
cc_264 N_A_XI20.X0_PGD N_B_c_568_n 0.00133285f
cc_265 N_A_c_343_n N_B_c_540_n 0.00124487f
cc_266 N_A_c_349_n N_B_c_540_n 0.00208788f
cc_267 N_A_c_361_n N_B_c_540_n 0.00263274f
cc_268 N_A_c_361_n N_Z_c_602_n 0.00109616f
cc_269 N_A_XI20.X0_PGD N_Z_c_606_n 7.88059e-19
cc_270 N_A_c_349_n N_Z_c_606_n 0.00136894f
cc_271 N_A_c_361_n N_Z_c_606_n 0.00142189f
cc_272 N_BI_c_456_p N_AI_XI19.X0_PGD 9.65637e-19
cc_273 N_BI_c_457_p N_AI_XI19.X0_PGD 0.00133285f
cc_274 N_BI_c_454_n N_AI_c_494_n 5.87796e-19
cc_275 N_BI_c_459_p N_AI_c_497_n 3.22026e-19
cc_276 N_BI_c_457_p N_AI_c_497_n 3.2351e-19
cc_277 N_BI_c_427_n N_AI_c_497_n 0.00274992f
cc_278 N_BI_c_455_n N_AI_c_497_n 2.49817e-19
cc_279 N_BI_c_459_p N_AI_c_506_n 3.26631e-19
cc_280 N_BI_c_457_p N_AI_c_506_n 0.00116273f
cc_281 N_BI_c_421_n N_B_c_538_n 6.8653e-19
cc_282 N_BI_c_423_n B 4.49325e-19
cc_283 N_BI_c_459_p N_B_c_562_n 6.00485e-19
cc_284 N_BI_c_457_p N_B_c_562_n 4.7755e-19
cc_285 N_BI_c_455_n N_B_c_562_n 3.12886e-19
cc_286 N_BI_c_438_n N_B_c_551_n 0.00178472f
cc_287 N_BI_c_459_p N_B_c_567_n 4.95293e-19
cc_288 N_BI_c_457_p N_B_c_567_n 0.00384234f
cc_289 N_BI_c_450_n N_B_c_567_n 6.17967e-19
cc_290 N_BI_c_438_n N_B_c_568_n 4.56568e-19
cc_291 N_BI_c_457_p N_B_c_568_n 7.16621e-19
cc_292 N_BI_c_450_n N_B_c_568_n 0.00243716f
cc_293 N_BI_c_438_n N_B_c_540_n 0.00166188f
cc_294 N_BI_c_455_n N_B_c_540_n 0.0081489f
cc_295 N_BI_c_430_n N_B_c_540_n 7.19198e-19
cc_296 N_BI_c_431_n N_B_c_540_n 8.87908e-19
cc_297 N_BI_c_455_n N_B_c_588_n 0.00345251f
cc_298 N_BI_c_482_p N_B_c_588_n 0.00190039f
cc_299 N_BI_c_430_n N_B_c_552_n 8.29167e-19
cc_300 N_BI_c_423_n N_B_c_550_n 0.00221197f
cc_301 N_BI_c_427_n N_B_c_550_n 0.0081489f
cc_302 N_BI_c_459_p N_Z_c_606_n 0.00181417f
cc_303 N_BI_c_438_n N_Z_c_606_n 0.00138952f
cc_304 N_BI_c_450_n N_Z_c_606_n 8.66889e-19
cc_305 N_BI_c_455_n N_Z_c_606_n 4.80971e-19
cc_306 N_AI_XI19.X0_PGD N_B_XI19.X0_CG 9.47088e-19
cc_307 N_AI_XI19.X0_PGD N_B_c_567_n 0.00133285f
cc_308 N_AI_XI19.X0_PGD N_Z_c_606_n 4.24145e-19
cc_309 N_B_c_562_n N_Z_c_606_n 0.00138952f
cc_310 N_B_c_551_n N_Z_c_606_n 0.00138952f
cc_311 N_B_c_567_n N_Z_c_606_n 8.66889e-19
cc_312 N_B_c_568_n N_Z_c_606_n 8.66889e-19
cc_313 N_B_c_540_n N_Z_c_606_n 0.0010571f
cc_314 N_B_c_588_n N_Z_c_606_n 0.00213616f
cc_315 N_B_c_552_n N_Z_c_606_n 0.00102447f
*
.ends
*
*
.subckt XNOR3_HPNW8 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XNOR3_N2
.ends
*
* File: G4_XOR2_N2.pex.netlist
* Created: Sun Apr 10 19:56:43 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XOR2_N2_VSS 2 5 9 12 14 16 32 33 42 43 45 54 59 63 66 71 76 81 86
+ 95 100 113 115 116 117 122 123 128 138 140 145 146 147 150
c98 148 0 6.15603e-19
c99 147 0 3.75522e-19
c100 146 0 4.28045e-19
c101 145 0 0.00386476f
c102 140 0 0.0021378f
c103 138 0 0.00844222f
c104 128 0 0.00339884f
c105 123 0 8.42592e-19
c106 122 0 0.00171246f
c107 117 0 8.20625e-19
c108 116 0 0.00418359f
c109 115 0 0.00524404f
c110 113 0 0.00159018f
c111 100 0 0.00404792f
c112 95 0 0.00404489f
c113 86 0 1.66825e-19
c114 81 0 0.00174451f
c115 76 0 6.28678e-19
c116 71 0 9.88359e-19
c117 66 0 0.00180488f
c118 63 0 0.00552459f
c119 59 0 0.00736499f
c120 54 0 0.00542864f
c121 45 0 1.03318e-19
c122 43 0 0.0342891f
c123 42 0 0.100068f
c124 33 0 0.0350852f
c125 32 0 0.0990727f
c126 14 0 0.00143442f
c127 9 0 0.269235f
c128 5 0 0.268907f
r129 145 150 0.326018
r130 144 145 4.58464
r131 140 144 0.655813
r132 139 148 0.494161
r133 138 150 0.326018
r134 138 139 13.0037
r135 134 148 0.128424
r136 129 147 0.494161
r137 128 148 0.494161
r138 128 129 7.46046
r139 124 147 0.128424
r140 122 147 0.494161
r141 122 123 4.37625
r142 118 146 0.0828784
r143 116 130 0.652036
r144 116 117 10.1279
r145 115 123 0.652036
r146 114 146 0.551426
r147 114 115 14.4208
r148 113 146 0.551426
r149 112 117 0.652036
r150 112 113 4.58464
r151 86 140 1.82344
r152 81 134 5.2515
r153 76 100 1.16709
r154 76 130 2.16729
r155 71 95 1.16709
r156 71 124 2.16729
r157 66 118 1.82344
r158 63 86 1.16709
r159 59 81 1.16709
r160 54 66 1.16709
r161 45 100 0.0476429
r162 43 45 1.45875
r163 42 46 0.652036
r164 42 45 1.45875
r165 39 43 0.652036
r166 35 95 0.0476429
r167 33 35 1.45875
r168 32 36 0.652036
r169 32 35 1.45875
r170 29 33 0.652036
r171 16 63 0.185659
r172 14 59 0.185659
r173 12 59 0.185659
r174 9 46 3.8511
r175 9 39 3.8511
r176 5 36 3.8511
r177 5 29 3.8511
r178 2 54 0.185659
.ends

.subckt PM_G4_XOR2_N2_VDD 3 6 8 11 14 16 32 42 43 54 59 63 66 68 69 70 73 75 76
+ 79 81 85 89 91 93 98 99 100 103 109 114
c99 114 0 0.00454282f
c100 109 0 0.00472544f
c101 101 0 8.79456e-19
c102 100 0 2.39889e-19
c103 99 0 4.52364e-19
c104 98 0 0.00483655f
c105 93 0 0.00147365f
c106 91 0 0.0130047f
c107 89 0 0.00227129f
c108 85 0 8.26969e-19
c109 81 0 0.00455615f
c110 79 0 0.00100252f
c111 76 0 8.63853e-19
c112 75 0 0.0057282f
c113 73 0 0.0019575f
c114 70 0 8.67926e-19
c115 69 0 0.00221146f
c116 68 0 0.00205498f
c117 66 0 0.00803904f
c118 63 0 0.00389115f
c119 59 0 0.00739215f
c120 54 0 0.00398638f
c121 43 0 0.0351228f
c122 42 0 0.100954f
c123 35 0 2.09107e-19
c124 33 0 0.035919f
c125 32 0 0.100953f
c126 14 0 0.00143442f
c127 11 0 0.269396f
c128 3 0 0.270542f
r129 98 103 0.349767
r130 97 98 4.58464
r131 93 103 0.306046
r132 93 95 1.82344
r133 92 101 0.494161
r134 91 97 0.652036
r135 91 92 13.0037
r136 87 101 0.128424
r137 87 89 5.2515
r138 85 114 1.16709
r139 83 85 2.16729
r140 82 100 0.494161
r141 81 101 0.494161
r142 81 82 7.46046
r143 79 109 1.16709
r144 77 100 0.128424
r145 77 79 2.16729
r146 75 83 0.652036
r147 75 76 10.1279
r148 71 99 0.0828784
r149 71 73 1.82344
r150 69 100 0.494161
r151 69 70 4.37625
r152 68 76 0.652036
r153 67 99 0.551426
r154 67 68 4.58464
r155 66 99 0.551426
r156 65 70 0.652036
r157 65 66 14.4208
r158 63 95 1.16709
r159 59 89 1.16709
r160 54 73 1.02121
r161 45 114 0.0476429
r162 43 45 1.45875
r163 42 46 0.652036
r164 42 45 1.45875
r165 39 43 0.652036
r166 35 109 0.0476429
r167 33 35 1.45875
r168 32 36 0.652036
r169 32 35 1.45875
r170 29 33 0.652036
r171 16 63 0.185659
r172 14 59 0.185659
r173 11 46 3.8511
r174 11 39 3.8511
r175 8 59 0.185659
r176 6 54 0.185659
r177 3 36 3.8511
r178 3 29 3.8511
.ends

.subckt PM_G4_XOR2_N2_A 2 4 7 10 21 24 28 39 48 51 54 57 62 67 72 77 85
c58 85 0 8.29046e-19
c59 77 0 0.00201173f
c60 72 0 0.00648506f
c61 67 0 0.00351476f
c62 62 0 0.00246599f
c63 57 0 0.00406665f
c64 54 0 7.62653e-19
c65 48 0 0.128037f
c66 43 0 0.0296312f
c67 39 0 2.38608e-19
c68 28 0 0.152668f
c69 24 0 9.84889e-20
c70 21 0 0.169628f
c71 18 0 0.126125f
c72 16 0 0.0247918f
c73 10 0 0.1218f
c74 7 0 0.324846f
c75 4 0 0.138512f
r76 81 85 0.653045
r77 62 77 1.16709
r78 62 85 4.9014
r79 57 72 1.16709
r80 57 81 9.00257
r81 54 67 1.16709
r82 51 54 0.0364688
r83 47 72 0.0238214
r84 47 48 2.334
r85 44 47 2.20433
r86 39 77 0.50025
r87 33 48 0.00605528
r88 31 44 0.00605528
r89 29 43 0.494161
r90 28 30 0.652036
r91 28 29 4.84305
r92 25 43 0.128424
r93 24 67 0.0476429
r94 22 24 0.326018
r95 22 24 0.1167
r96 21 43 0.494161
r97 21 24 6.7686
r98 18 67 0.357321
r99 16 24 0.326018
r100 16 18 0.40845
r101 10 39 3.3843
r102 7 33 3.8511
r103 7 31 3.8511
r104 7 30 3.8511
r105 4 25 3.8511
r106 2 18 3.44265
.ends

.subckt PM_G4_XOR2_N2_NET1 2 4 7 10 30 31 35 41 44 49 58 76
c37 76 0 3.4517e-19
c38 58 0 0.00413905f
c39 49 0 0.00667491f
c40 44 0 0.00198364f
c41 41 0 0.00539823f
c42 35 0 0.103124f
c43 31 0 0.125482f
c44 30 0 9.62407e-20
c45 10 0 0.214624f
c46 7 0 0.384182f
c47 4 0 0.00143442f
r48 72 76 0.655813
r49 49 58 1.16709
r50 49 76 12.1076
r51 44 72 2.41736
r52 41 44 1.16709
r53 33 35 1.70187
r54 30 58 0.0238214
r55 30 31 2.20433
r56 27 30 2.334
r57 25 35 0.17282
r58 24 31 0.00605528
r59 21 33 0.17282
r60 18 27 0.00605528
r61 10 21 6.36015
r62 7 25 6.01005
r63 7 24 3.8511
r64 7 18 3.8511
r65 4 41 0.185659
r66 2 41 0.185659
.ends

.subckt PM_G4_XOR2_N2_NET2 2 4 6 9 21 22 33 39 42 47 56 74
c44 74 0 3.04338e-19
c45 56 0 0.00509819f
c46 47 0 0.00799947f
c47 42 0 0.00221316f
c48 39 0 0.00534974f
c49 33 0 0.129063f
c50 22 0 0.0345383f
c51 21 0 0.17396f
c52 9 0 0.466016f
c53 6 0 0.135514f
c54 4 0 0.00143442f
r55 70 74 0.660011
r56 47 56 1.16709
r57 47 74 11.3611
r58 42 70 2.37568
r59 39 42 1.16709
r60 32 56 0.0238214
r61 32 33 2.26917
r62 29 32 2.26917
r63 26 33 0.00605528
r64 24 29 0.00605528
r65 21 23 0.652036
r66 21 22 4.84305
r67 18 22 0.652036
r68 9 26 3.8511
r69 9 24 3.8511
r70 9 23 8.7525
r71 6 18 3.8511
r72 4 39 0.185659
r73 2 39 0.185659
.ends

.subckt PM_G4_XOR2_N2_B 2 4 7 10 19 20 28 31 35 45 52 55
c33 55 0 0.0280361f
c34 52 0 0.00155244f
c35 45 0 0.13326f
c36 35 0 0.154246f
c37 31 0 9.67975e-20
c38 28 0 0.117533f
c39 20 0 0.0348105f
c40 19 0 0.169544f
c41 10 0 0.209756f
c42 7 0 0.32787f
c43 4 0 0.134866f
c44 2 0 0.146861f
r45 49 55 1.16709
r46 49 52 0.0364688
r47 43 45 4.53833
r48 38 45 0.00605528
r49 35 47 1.87725
r50 33 47 0.527901
r51 32 43 0.00605528
r52 31 55 0.181909
r53 29 55 0.494161
r54 29 31 0.1167
r55 28 47 0.333556
r56 28 31 4.72635
r57 23 55 0.128424
r58 23 55 0.40845
r59 22 55 0.181909
r60 20 22 6.7686
r61 19 55 0.494161
r62 19 22 0.1167
r63 16 20 0.652036
r64 10 35 6.3018
r65 7 38 3.8511
r66 7 33 4.14285
r67 7 32 3.8511
r68 4 55 3.7344
r69 2 16 4.14285
.ends

.subckt PM_G4_XOR2_N2_Z 2 4 6 8 23 27 30 33
c29 30 0 0.00340522f
c30 27 0 0.00725263f
c31 23 0 0.0052085f
c32 8 0 0.00143442f
c33 6 0 0.00143442f
r34 33 35 3.83443
r35 30 33 6.00171
r36 27 35 1.16709
r37 23 30 1.16709
r38 8 27 0.185659
r39 6 23 0.185659
r40 4 27 0.185659
r41 2 23 0.185659
.ends

.subckt G4_XOR2_N2  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI14.X0 N_NET1_XI14.X0_D N_VDD_XI14.X0_PGD N_B_XI14.X0_CG N_VDD_XI14.X0_PGD
+ N_VSS_XI14.X0_S TIGFET_HPNW8
XI4.X0 N_NET2_XI4.X0_D N_VSS_XI4.X0_PGD N_A_XI4.X0_CG N_VSS_XI4.X0_PGD
+ N_VDD_XI4.X0_S TIGFET_HPNW8
XI12.X0 N_NET1_XI12.X0_D N_VSS_XI12.X0_PGD N_B_XI12.X0_CG N_VSS_XI12.X0_PGD
+ N_VDD_XI12.X0_S TIGFET_HPNW8
XI0.X0 N_NET2_XI0.X0_D N_VDD_XI0.X0_PGD N_A_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW8
XI15.X0 N_Z_XI15.X0_D N_B_XI15.X0_PGD N_NET2_XI15.X0_CG N_B_XI15.X0_PGD
+ N_VDD_XI15.X0_S TIGFET_HPNW8
XI6.X0 N_Z_XI6.X0_D N_A_XI6.X0_PGD N_B_XI6.X0_CG N_A_XI6.X0_PGD N_VSS_XI6.X0_S
+ TIGFET_HPNW8
XI13.X0 N_Z_XI13.X0_D N_NET1_XI13.X0_PGD N_A_XI13.X0_CG N_NET1_XI13.X0_PGD
+ N_VDD_XI13.X0_S TIGFET_HPNW8
XI2.X0 N_Z_XI2.X0_D N_NET2_XI2.X0_PGD N_NET1_XI2.X0_CG N_NET2_XI2.X0_PGD
+ N_VSS_XI2.X0_S TIGFET_HPNW8
*
x_PM_G4_XOR2_N2_VSS N_VSS_XI14.X0_S N_VSS_XI4.X0_PGD N_VSS_XI12.X0_PGD
+ N_VSS_XI0.X0_S N_VSS_XI6.X0_S N_VSS_XI2.X0_S N_VSS_c_5_p N_VSS_c_22_p
+ N_VSS_c_37_p N_VSS_c_4_p N_VSS_c_84_p N_VSS_c_7_p N_VSS_c_6_p N_VSS_c_91_p
+ N_VSS_c_8_p N_VSS_c_13_p N_VSS_c_29_p N_VSS_c_35_p N_VSS_c_39_p N_VSS_c_14_p
+ N_VSS_c_32_p N_VSS_c_9_p N_VSS_c_10_p N_VSS_c_18_p N_VSS_c_19_p N_VSS_c_25_p
+ N_VSS_c_28_p N_VSS_c_26_p N_VSS_c_55_p N_VSS_c_40_p N_VSS_c_77_p N_VSS_c_11_p
+ N_VSS_c_27_p VSS PM_G4_XOR2_N2_VSS
x_PM_G4_XOR2_N2_VDD N_VDD_XI14.X0_PGD N_VDD_XI4.X0_S N_VDD_XI12.X0_S
+ N_VDD_XI0.X0_PGD N_VDD_XI15.X0_S N_VDD_XI13.X0_S N_VDD_c_102_n N_VDD_c_149_p
+ N_VDD_c_103_n N_VDD_c_175_p N_VDD_c_104_n N_VDD_c_189_p N_VDD_c_105_n
+ N_VDD_c_110_n N_VDD_c_114_n N_VDD_c_117_n N_VDD_c_118_n N_VDD_c_119_n
+ N_VDD_c_126_n N_VDD_c_127_n N_VDD_c_128_n N_VDD_c_132_n N_VDD_c_135_n
+ N_VDD_c_154_p N_VDD_c_137_n N_VDD_c_162_p N_VDD_c_139_n N_VDD_c_140_n VDD
+ N_VDD_c_141_n N_VDD_c_143_n PM_G4_XOR2_N2_VDD
x_PM_G4_XOR2_N2_A N_A_XI4.X0_CG N_A_XI0.X0_CG N_A_XI6.X0_PGD N_A_XI13.X0_CG
+ N_A_c_198_n N_A_c_200_n N_A_c_201_n N_A_c_230_p N_A_c_216_n A N_A_c_202_n
+ N_A_c_204_n N_A_c_208_n N_A_c_209_n N_A_c_225_n N_A_c_229_p N_A_c_211_n
+ PM_G4_XOR2_N2_A
x_PM_G4_XOR2_N2_NET1 N_NET1_XI14.X0_D N_NET1_XI12.X0_D N_NET1_XI13.X0_PGD
+ N_NET1_XI2.X0_CG N_NET1_c_279_n N_NET1_c_263_n N_NET1_c_284_p N_NET1_c_256_n
+ N_NET1_c_257_n N_NET1_c_259_n N_NET1_c_273_n N_NET1_c_261_n PM_G4_XOR2_N2_NET1
x_PM_G4_XOR2_N2_NET2 N_NET2_XI4.X0_D N_NET2_XI0.X0_D N_NET2_XI15.X0_CG
+ N_NET2_XI2.X0_PGD N_NET2_c_315_n N_NET2_c_331_p N_NET2_c_316_n N_NET2_c_293_n
+ N_NET2_c_295_n N_NET2_c_299_n N_NET2_c_321_n N_NET2_c_303_n PM_G4_XOR2_N2_NET2
x_PM_G4_XOR2_N2_B N_B_XI14.X0_CG N_B_XI12.X0_CG N_B_XI15.X0_PGD N_B_XI6.X0_CG
+ N_B_c_338_n N_B_c_356_n N_B_c_340_n N_B_c_341_n N_B_c_358_n N_B_c_342_n B
+ N_B_c_345_n PM_G4_XOR2_N2_B
x_PM_G4_XOR2_N2_Z N_Z_XI15.X0_D N_Z_XI6.X0_D N_Z_XI13.X0_D N_Z_XI2.X0_D
+ N_Z_c_379_n N_Z_c_370_n N_Z_c_374_n Z PM_G4_XOR2_N2_Z
cc_1 N_VSS_XI4.X0_PGD N_VDD_XI14.X0_PGD 3.09777e-19
cc_2 N_VSS_XI12.X0_PGD N_VDD_XI14.X0_PGD 0.0019593f
cc_3 N_VSS_XI4.X0_PGD N_VDD_XI0.X0_PGD 0.0019696f
cc_4 N_VSS_c_4_p N_VDD_c_102_n 0.0019593f
cc_5 N_VSS_c_5_p N_VDD_c_103_n 0.0019696f
cc_6 N_VSS_c_6_p N_VDD_c_104_n 3.3848e-19
cc_7 N_VSS_c_7_p N_VDD_c_105_n 9.5668e-19
cc_8 N_VSS_c_8_p N_VDD_c_105_n 0.00165395f
cc_9 N_VSS_c_9_p N_VDD_c_105_n 0.00337557f
cc_10 N_VSS_c_10_p N_VDD_c_105_n 0.00738982f
cc_11 N_VSS_c_11_p N_VDD_c_105_n 9.16632e-19
cc_12 N_VSS_XI4.X0_PGD N_VDD_c_110_n 2.76462e-19
cc_13 N_VSS_c_13_p N_VDD_c_110_n 4.35319e-19
cc_14 N_VSS_c_14_p N_VDD_c_110_n 3.66936e-19
cc_15 N_VSS_c_10_p N_VDD_c_110_n 0.00312786f
cc_16 N_VSS_c_7_p N_VDD_c_114_n 3.4118e-19
cc_17 N_VSS_c_8_p N_VDD_c_114_n 4.19648e-19
cc_18 N_VSS_c_18_p N_VDD_c_114_n 0.0035394f
cc_19 N_VSS_c_19_p N_VDD_c_117_n 0.00106066f
cc_20 N_VSS_c_8_p N_VDD_c_118_n 5.20373e-19
cc_21 N_VSS_c_5_p N_VDD_c_119_n 3.9313e-19
cc_22 N_VSS_c_22_p N_VDD_c_119_n 3.9313e-19
cc_23 N_VSS_c_13_p N_VDD_c_119_n 0.00141228f
cc_24 N_VSS_c_14_p N_VDD_c_119_n 0.00114511f
cc_25 N_VSS_c_25_p N_VDD_c_119_n 0.00345257f
cc_26 N_VSS_c_26_p N_VDD_c_119_n 0.00601358f
cc_27 N_VSS_c_27_p N_VDD_c_119_n 7.74609e-19
cc_28 N_VSS_c_28_p N_VDD_c_126_n 0.00107662f
cc_29 N_VSS_c_29_p N_VDD_c_127_n 9.53862e-19
cc_30 N_VSS_c_4_p N_VDD_c_128_n 3.9313e-19
cc_31 N_VSS_c_29_p N_VDD_c_128_n 0.00161703f
cc_32 N_VSS_c_32_p N_VDD_c_128_n 2.26455e-19
cc_33 N_VSS_c_18_p N_VDD_c_128_n 0.0060445f
cc_34 N_VSS_c_13_p N_VDD_c_132_n 9.25722e-19
cc_35 N_VSS_c_35_p N_VDD_c_132_n 9.24903e-19
cc_36 N_VSS_c_14_p N_VDD_c_132_n 3.99794e-19
cc_37 N_VSS_c_37_p N_VDD_c_135_n 2.36788e-19
cc_38 N_VSS_c_29_p N_VDD_c_135_n 0.00251632f
cc_39 N_VSS_c_39_p N_VDD_c_137_n 2.22977e-19
cc_40 N_VSS_c_40_p N_VDD_c_137_n 0.00110879f
cc_41 N_VSS_c_10_p N_VDD_c_139_n 0.0010705f
cc_42 N_VSS_c_18_p N_VDD_c_140_n 0.00108916f
cc_43 N_VSS_c_29_p N_VDD_c_141_n 3.48267e-19
cc_44 N_VSS_c_32_p N_VDD_c_141_n 6.46219e-19
cc_45 N_VSS_c_13_p N_VDD_c_143_n 3.48267e-19
cc_46 N_VSS_c_14_p N_VDD_c_143_n 6.489e-19
cc_47 N_VSS_XI4.X0_PGD N_A_c_198_n 4.04227e-19
cc_48 N_VSS_XI12.X0_PGD N_A_c_198_n 2.49256e-19
cc_49 N_VSS_c_14_p N_A_c_200_n 9.46927e-19
cc_50 N_VSS_XI12.X0_PGD N_A_c_201_n 2.49256e-19
cc_51 N_VSS_c_13_p N_A_c_202_n 3.33636e-19
cc_52 N_VSS_c_14_p N_A_c_202_n 3.2351e-19
cc_53 N_VSS_c_35_p N_A_c_204_n 0.00580642f
cc_54 N_VSS_c_10_p N_A_c_204_n 7.28437e-19
cc_55 N_VSS_c_55_p N_A_c_204_n 0.00192457f
cc_56 N_VSS_c_40_p N_A_c_204_n 3.96468e-19
cc_57 N_VSS_c_55_p N_A_c_208_n 6.42713e-19
cc_58 N_VSS_c_13_p N_A_c_209_n 3.2351e-19
cc_59 N_VSS_c_14_p N_A_c_209_n 2.68747e-19
cc_60 N_VSS_c_55_p N_A_c_211_n 4.97622e-19
cc_61 N_VSS_c_7_p N_NET1_c_256_n 3.43419e-19
cc_62 N_VSS_c_8_p N_NET1_c_257_n 0.00115894f
cc_63 N_VSS_c_18_p N_NET1_c_257_n 2.79692e-19
cc_64 N_VSS_c_29_p N_NET1_c_259_n 0.00143375f
cc_65 N_VSS_c_35_p N_NET1_c_259_n 2.33463e-19
cc_66 N_VSS_c_9_p N_NET1_c_261_n 4.42442e-19
cc_67 N_VSS_c_18_p N_NET1_c_261_n 4.73555e-19
cc_68 N_VSS_c_6_p N_NET2_c_293_n 3.43419e-19
cc_69 N_VSS_c_35_p N_NET2_c_293_n 3.48267e-19
cc_70 N_VSS_c_6_p N_NET2_c_295_n 3.48267e-19
cc_71 N_VSS_c_35_p N_NET2_c_295_n 0.00163864f
cc_72 N_VSS_c_10_p N_NET2_c_295_n 6.00032e-19
cc_73 N_VSS_c_26_p N_NET2_c_295_n 2.79074e-19
cc_74 N_VSS_c_35_p N_NET2_c_299_n 0.00185959f
cc_75 N_VSS_c_26_p N_NET2_c_299_n 0.00111941f
cc_76 N_VSS_c_55_p N_NET2_c_299_n 0.0051115f
cc_77 N_VSS_c_77_p N_NET2_c_299_n 0.00115623f
cc_78 N_VSS_c_13_p N_NET2_c_303_n 5.67902e-19
cc_79 N_VSS_c_26_p N_NET2_c_303_n 4.76092e-19
cc_80 N_VSS_XI12.X0_PGD N_B_XI15.X0_PGD 0.00190378f
cc_81 N_VSS_XI4.X0_PGD N_B_c_338_n 2.59761e-19
cc_82 N_VSS_XI12.X0_PGD N_B_c_338_n 4.04459e-19
cc_83 N_VSS_XI12.X0_PGD N_B_c_340_n 4.08222e-19
cc_84 N_VSS_c_84_p N_B_c_341_n 8.74538e-19
cc_85 N_VSS_c_37_p N_B_c_342_n 0.00168656f
cc_86 N_VSS_c_29_p B 3.14335e-19
cc_87 N_VSS_c_32_p B 3.07907e-19
cc_88 N_VSS_c_29_p N_B_c_345_n 3.07907e-19
cc_89 N_VSS_c_32_p N_B_c_345_n 2.38856e-19
cc_90 N_VSS_c_6_p N_Z_c_370_n 3.43419e-19
cc_91 N_VSS_c_91_p N_Z_c_370_n 3.43419e-19
cc_92 N_VSS_c_35_p N_Z_c_370_n 3.48267e-19
cc_93 N_VSS_c_39_p N_Z_c_370_n 3.48267e-19
cc_94 N_VSS_c_6_p N_Z_c_374_n 3.48267e-19
cc_95 N_VSS_c_91_p N_Z_c_374_n 3.48267e-19
cc_96 N_VSS_c_35_p N_Z_c_374_n 4.84964e-19
cc_97 N_VSS_c_39_p N_Z_c_374_n 5.71987e-19
cc_98 N_VSS_c_55_p N_Z_c_374_n 3.24575e-19
cc_99 N_VDD_XI0.X0_PGD N_A_XI6.X0_PGD 0.00170367f
cc_100 N_VDD_XI14.X0_PGD N_A_c_198_n 2.49256e-19
cc_101 N_VDD_XI0.X0_PGD N_A_c_198_n 4.07423e-19
cc_102 N_VDD_XI0.X0_PGD N_A_c_201_n 4.08222e-19
cc_103 N_VDD_c_149_p N_A_c_216_n 0.00170367f
cc_104 N_VDD_c_105_n N_A_c_202_n 5.04211e-19
cc_105 N_VDD_c_127_n N_A_c_202_n 2.0061e-19
cc_106 N_VDD_c_132_n N_A_c_204_n 4.55539e-19
cc_107 N_VDD_c_143_n N_A_c_204_n 3.5189e-19
cc_108 N_VDD_c_154_p N_A_c_208_n 6.92642e-19
cc_109 N_VDD_c_105_n N_A_c_209_n 5.74039e-19
cc_110 N_VDD_c_127_n N_A_c_209_n 2.00694e-19
cc_111 N_VDD_c_141_n N_A_c_209_n 2.58157e-19
cc_112 N_VDD_c_132_n N_A_c_225_n 4.08069e-19
cc_113 N_VDD_c_143_n N_A_c_225_n 6.61916e-19
cc_114 N_VDD_c_154_p N_A_c_211_n 8.87092e-19
cc_115 N_VDD_c_154_p N_NET1_c_263_n 8.59992e-19
cc_116 N_VDD_c_162_p N_NET1_c_263_n 2.76493e-19
cc_117 N_VDD_c_104_n N_NET1_c_256_n 3.43419e-19
cc_118 N_VDD_c_135_n N_NET1_c_256_n 3.48267e-19
cc_119 N_VDD_c_104_n N_NET1_c_257_n 3.48267e-19
cc_120 N_VDD_c_128_n N_NET1_c_257_n 4.34701e-19
cc_121 N_VDD_c_135_n N_NET1_c_257_n 0.00119216f
cc_122 N_VDD_c_135_n N_NET1_c_259_n 0.00121188f
cc_123 N_VDD_c_154_p N_NET1_c_259_n 0.00357992f
cc_124 N_VDD_c_162_p N_NET1_c_259_n 8.17443e-19
cc_125 N_VDD_c_135_n N_NET1_c_273_n 2.78343e-19
cc_126 N_VDD_c_154_p N_NET1_c_273_n 2.67643e-19
cc_127 N_VDD_c_162_p N_NET1_c_273_n 3.70842e-19
cc_128 N_VDD_c_127_n N_NET1_c_261_n 2.94681e-19
cc_129 N_VDD_c_175_p N_NET2_c_293_n 3.67949e-19
cc_130 N_VDD_c_118_n N_NET2_c_293_n 3.72199e-19
cc_131 N_VDD_c_175_p N_NET2_c_295_n 3.9802e-19
cc_132 N_VDD_c_118_n N_NET2_c_295_n 5.226e-19
cc_133 N_VDD_c_119_n N_NET2_c_295_n 4.34701e-19
cc_134 N_VDD_c_132_n N_NET2_c_299_n 2.89449e-19
cc_135 N_VDD_c_105_n N_B_XI14.X0_CG 3.86879e-19
cc_136 N_VDD_XI14.X0_PGD N_B_c_338_n 4.0747e-19
cc_137 N_VDD_XI0.X0_PGD N_B_c_338_n 2.59761e-19
cc_138 N_VDD_XI0.X0_PGD N_B_c_340_n 2.59761e-19
cc_139 N_VDD_c_135_n N_B_c_342_n 2.45557e-19
cc_140 N_VDD_c_154_p N_B_c_342_n 0.00104936f
cc_141 N_VDD_c_143_n N_B_c_345_n 3.88194e-19
cc_142 N_VDD_c_104_n N_Z_c_379_n 3.43419e-19
cc_143 N_VDD_c_189_p N_Z_c_379_n 3.43419e-19
cc_144 N_VDD_c_135_n N_Z_c_379_n 3.48267e-19
cc_145 N_VDD_c_154_p N_Z_c_379_n 3.4118e-19
cc_146 N_VDD_c_137_n N_Z_c_379_n 3.72199e-19
cc_147 N_VDD_c_104_n N_Z_c_374_n 3.48267e-19
cc_148 N_VDD_c_189_p N_Z_c_374_n 3.48267e-19
cc_149 N_VDD_c_135_n N_Z_c_374_n 7.9714e-19
cc_150 N_VDD_c_154_p N_Z_c_374_n 6.28755e-19
cc_151 N_VDD_c_137_n N_Z_c_374_n 8.5731e-19
cc_152 N_A_XI13.X0_CG N_NET1_XI13.X0_PGD 9.16948e-19
cc_153 N_A_c_229_p N_NET1_XI13.X0_PGD 5.82245e-19
cc_154 N_A_c_230_p N_NET1_c_279_n 8.72031e-19
cc_155 N_A_c_208_n N_NET1_c_259_n 0.00253116f
cc_156 N_A_c_211_n N_NET1_c_259_n 6.96104e-19
cc_157 N_A_c_229_p N_NET1_c_273_n 2.38856e-19
cc_158 N_A_XI13.X0_CG N_NET2_XI15.X0_CG 2.29068e-19
cc_159 N_A_XI6.X0_PGD N_NET2_XI2.X0_PGD 0.00174971f
cc_160 N_A_c_201_n N_NET2_XI2.X0_PGD 3.14428e-19
cc_161 N_A_c_229_p N_NET2_XI2.X0_PGD 3.71891e-19
cc_162 N_A_XI6.X0_PGD N_NET2_c_315_n 4.63684e-19
cc_163 N_A_c_216_n N_NET2_c_316_n 0.00174971f
cc_164 N_A_c_198_n N_NET2_c_293_n 5.99889e-19
cc_165 N_A_c_204_n N_NET2_c_299_n 0.0021219f
cc_166 N_A_c_208_n N_NET2_c_299_n 0.00109012f
cc_167 N_A_c_225_n N_NET2_c_299_n 3.44698e-19
cc_168 N_A_c_230_p N_NET2_c_321_n 4.27572e-19
cc_169 N_A_c_204_n N_NET2_c_321_n 3.44698e-19
cc_170 N_A_c_225_n N_NET2_c_321_n 6.78604e-19
cc_171 N_A_c_201_n N_B_XI6.X0_CG 0.003858f
cc_172 N_A_c_198_n N_B_c_338_n 0.00631299f
cc_173 N_A_c_209_n N_B_c_356_n 8.20069e-19
cc_174 N_A_c_201_n N_B_c_340_n 0.00464284f
cc_175 N_A_c_201_n N_B_c_358_n 0.00220484f
cc_176 N_A_c_198_n N_B_c_345_n 8.92181e-19
cc_177 N_A_c_204_n N_Z_c_374_n 0.00336431f
cc_178 N_A_c_208_n N_Z_c_374_n 0.00291096f
cc_179 N_A_c_229_p N_Z_c_374_n 9.75659e-19
cc_180 N_NET1_XI13.X0_PGD N_NET2_XI15.X0_CG 2.3921e-19
cc_181 N_NET1_c_284_p N_NET2_XI2.X0_PGD 0.00790765f
cc_182 N_NET1_XI13.X0_PGD N_NET2_c_315_n 0.00383f
cc_183 N_NET1_c_256_n N_NET2_c_293_n 2.51993e-19
cc_184 N_NET1_XI13.X0_PGD N_B_XI15.X0_PGD 0.00215865f
cc_185 N_NET1_XI2.X0_CG N_B_XI6.X0_CG 2.58346e-19
cc_186 N_NET1_c_256_n N_B_c_338_n 5.53604e-19
cc_187 N_NET1_c_284_p N_B_c_358_n 2.58346e-19
cc_188 N_NET1_c_263_n N_B_c_342_n 0.00193302f
cc_189 N_NET1_c_259_n N_Z_c_374_n 2.36895e-19
cc_190 N_NET2_XI15.X0_CG N_B_XI15.X0_PGD 0.00204226f
cc_191 N_NET2_c_315_n N_B_XI15.X0_PGD 0.00161654f
cc_192 N_NET2_XI2.X0_PGD N_B_c_358_n 0.00351134f
cc_193 N_NET2_c_331_p N_B_c_358_n 0.00396313f
cc_194 N_NET2_c_315_n N_Z_c_379_n 7.46018e-19
cc_195 N_NET2_c_315_n N_Z_c_370_n 2.51166e-19
cc_196 N_NET2_XI2.X0_PGD N_Z_c_374_n 0.0012102f
cc_197 N_NET2_c_315_n N_Z_c_374_n 2.5304e-19
cc_198 N_NET2_c_299_n N_Z_c_374_n 3.59687e-19
cc_199 N_B_c_358_n N_Z_c_374_n 0.00106974f
*
.ends
*
*
.subckt XOR2_HPNW8 A B Y VDD VSS
xgate (VSS VDD A B Y) G4_XOR2_N2
.ends
*
* File: G5_XOR3_N2.pex.netlist
* Created: Thu Mar 31 11:38:36 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XOR3_N2_VDD 2 5 9 12 14 17 34 35 44 45 47 54 55 65 69 74 77 79 80
+ 81 84 86 90 93 96 98 102 104 108 112 114 116 118 119 125 134 139 Vss
c115 139 Vss 0.00504502f
c116 134 Vss 0.00507145f
c117 125 Vss 0.00564924f
c118 119 Vss 2.39889e-19
c119 118 Vss 4.91626e-19
c120 117 Vss 5.50975e-19
c121 114 Vss 4.52364e-19
c122 112 Vss 0.00169191f
c123 108 Vss 0.00106552f
c124 104 Vss 0.00630988f
c125 102 Vss 0.00113412f
c126 98 Vss 0.00579331f
c127 96 Vss 0.00150773f
c128 93 Vss 0.00256047f
c129 90 Vss 0.00487749f
c130 86 Vss 0.00657827f
c131 84 Vss 0.00152345f
c132 81 Vss 8.67722e-19
c133 80 Vss 0.00905163f
c134 79 Vss 0.0103203f
c135 77 Vss 0.00223293f
c136 74 Vss 0.00377995f
c137 69 Vss 0.00394389f
c138 65 Vss 0.00382792f
c139 55 Vss 0.035607f
c140 54 Vss 0.100823f
c141 47 Vss 8.75732e-20
c142 45 Vss 0.0356105f
c143 44 Vss 0.101295f
c144 35 Vss 0.0346386f
c145 34 Vss 0.0990802f
c146 17 Vss 0.269219f
c147 9 Vss 0.270254f
c148 5 Vss 0.27424f
r149 110 112 5.2515
r150 108 139 1.16709
r151 106 108 2.16729
r152 105 119 0.494161
r153 104 110 0.652036
r154 104 105 7.46046
r155 102 134 1.16709
r156 100 119 0.128424
r157 100 102 2.16729
r158 99 118 0.494161
r159 98 106 0.652036
r160 98 99 10.3363
r161 94 117 0.0828784
r162 94 96 2.00578
r163 93 118 0.128424
r164 92 117 0.551426
r165 92 93 4.58464
r166 90 125 1.16709
r167 88 117 0.551426
r168 88 90 6.79361
r169 87 116 0.326018
r170 86 118 0.494161
r171 86 87 10.1279
r172 82 114 0.0828784
r173 82 84 1.82344
r174 80 119 0.494161
r175 80 81 15.8795
r176 79 116 0.326018
r177 78 114 0.551426
r178 78 79 15.6295
r179 77 114 0.551426
r180 76 81 0.652036
r181 76 77 4.58464
r182 74 112 1.16709
r183 69 96 1.16709
r184 65 84 1.16709
r185 57 139 0.0476429
r186 55 57 1.45875
r187 54 58 0.652036
r188 54 57 1.45875
r189 51 55 0.652036
r190 47 134 0.0476429
r191 45 47 1.45875
r192 44 48 0.652036
r193 44 47 1.45875
r194 41 45 0.652036
r195 37 125 0.238214
r196 35 37 1.45875
r197 34 38 0.652036
r198 34 37 1.45875
r199 31 35 0.652036
r200 17 58 3.8511
r201 17 51 3.8511
r202 14 74 0.185659
r203 12 69 0.185659
r204 9 48 3.8511
r205 9 41 3.8511
r206 5 38 3.8511
r207 5 31 3.8511
r208 2 65 0.185659
.ends

.subckt PM_G5_XOR3_N2_C 2 4 6 8 17 20 23 32 37 40 43 47 52 57 84 92 98 Vss
c55 98 Vss 3.07681e-19
c56 92 Vss 0.00543335f
c57 84 Vss 0.00807877f
c58 57 Vss 0.00478462f
c59 52 Vss 0.00202371f
c60 47 Vss 0.00149319f
c61 43 Vss 5.64514e-19
c62 40 Vss 6.40888e-19
c63 37 Vss 0.00399277f
c64 32 Vss 0.00492048f
c65 23 Vss 2.41681e-19
c66 20 Vss 0.221837f
c67 17 Vss 0.126125f
c68 15 Vss 0.0247918f
c69 4 Vss 0.133869f
r70 93 98 0.441572
r71 92 94 0.655813
r72 92 93 9.04425
r73 88 98 0.174814
r74 84 98 0.441572
r75 52 94 2.45904
r76 47 88 2.45904
r77 43 57 1.16709
r78 43 84 22.1365
r79 40 43 0.0416786
r80 37 52 1.16709
r81 32 47 1.16709
r82 23 57 0.0476429
r83 21 23 0.326018
r84 21 23 0.1167
r85 20 24 0.652036
r86 20 23 6.7686
r87 17 57 0.357321
r88 15 23 0.326018
r89 15 17 0.40845
r90 8 37 0.185659
r91 6 32 0.185659
r92 4 24 3.8511
r93 2 17 3.44265
.ends

.subckt PM_G5_XOR3_N2_VSS 3 6 8 11 15 18 34 37 44 45 54 55 57 66 70 73 78 83 88
+ 93 98 107 112 121 123 124 125 130 131 136 142 148 152 153 154 156 Vss
c125 154 Vss 3.75522e-19
c126 153 Vss 3.88979e-19
c127 152 Vss 4.4306e-19
c128 148 Vss 4.18562e-19
c129 142 Vss 0.00192878f
c130 136 Vss 0.00349848f
c131 131 Vss 8.4146e-19
c132 130 Vss 0.00631713f
c133 125 Vss 8.38522e-19
c134 124 Vss 0.00567123f
c135 123 Vss 0.00379369f
c136 121 Vss 0.00292495f
c137 112 Vss 0.00392167f
c138 107 Vss 0.00408825f
c139 98 Vss 0.00496033f
c140 93 Vss 0.00183916f
c141 88 Vss 6.78589e-19
c142 83 Vss 8.07476e-19
c143 78 Vss 0.00294517f
c144 73 Vss 0.00293431f
c145 70 Vss 0.00527641f
c146 66 Vss 0.00738472f
c147 57 Vss 1.05421e-19
c148 55 Vss 0.0347733f
c149 54 Vss 0.0996929f
c150 45 Vss 0.035088f
c151 44 Vss 0.0994129f
c152 37 Vss 6.29003e-20
c153 35 Vss 0.0348882f
c154 34 Vss 0.100326f
c155 15 Vss 0.270318f
c156 11 Vss 0.269056f
c157 8 Vss 0.00143442f
c158 3 Vss 0.275257f
r159 148 156 0.326018
r160 143 154 0.494161
r161 142 156 0.326018
r162 142 143 7.46046
r163 138 154 0.128424
r164 137 153 0.494161
r165 136 144 0.652036
r166 136 137 7.46046
r167 132 153 0.128424
r168 130 154 0.494161
r169 130 131 15.8795
r170 126 152 0.0828784
r171 124 153 0.494161
r172 124 125 13.0037
r173 123 131 0.652036
r174 122 152 0.551426
r175 122 123 12.0451
r176 121 152 0.551426
r177 120 125 0.652036
r178 120 121 8.169
r179 93 148 5.2515
r180 88 112 1.16709
r181 88 144 2.16729
r182 83 107 1.16709
r183 83 138 2.16729
r184 78 132 5.2515
r185 73 98 1.16709
r186 73 126 4.33978
r187 70 93 1.16709
r188 66 78 1.16709
r189 57 112 0.0476429
r190 55 57 1.45875
r191 54 58 0.652036
r192 54 57 1.45875
r193 51 55 0.652036
r194 47 107 0.0476429
r195 45 47 1.45875
r196 44 48 0.652036
r197 44 47 1.45875
r198 41 45 0.652036
r199 37 98 0.238214
r200 35 37 1.45875
r201 34 38 0.652036
r202 34 37 1.45875
r203 31 35 0.652036
r204 18 70 0.185659
r205 15 58 3.8511
r206 15 51 3.8511
r207 11 48 3.8511
r208 11 41 3.8511
r209 8 66 0.185659
r210 6 66 0.185659
r211 3 38 3.8511
r212 3 31 3.8511
.ends

.subckt PM_G5_XOR3_N2_CI 2 4 6 8 23 26 31 34 39 44 79 80 82 84 89 Vss
c55 95 Vss 8.69704e-20
c56 89 Vss 0.00497463f
c57 84 Vss 1.28221e-19
c58 83 Vss 1.74838e-19
c59 82 Vss 0.0011265f
c60 80 Vss 4.20409e-19
c61 79 Vss 0.00494114f
c62 44 Vss 0.00209131f
c63 39 Vss 0.00145787f
c64 34 Vss 0.00360912f
c65 31 Vss 0.00501643f
c66 26 Vss 0.00386883f
c67 23 Vss 0.00546777f
c68 4 Vss 0.00143442f
r69 90 95 0.494161
r70 89 91 0.652036
r71 89 90 10.3363
r72 85 95 0.128424
r73 83 95 0.494161
r74 83 84 1.70882
r75 82 84 0.652036
r76 81 82 4.75136
r77 79 81 0.652036
r78 79 80 18.9638
r79 75 80 0.652036
r80 44 91 2.58407
r81 39 85 2.58407
r82 34 75 7.71054
r83 31 44 1.16709
r84 26 39 1.16709
r85 23 34 1.16709
r86 8 31 0.185659
r87 6 26 0.185659
r88 4 23 0.185659
r89 2 23 0.185659
.ends

.subckt PM_G5_XOR3_N2_A 2 4 7 11 24 44 45 49 51 54 56 57 60 65 66 69 74 Vss
c72 74 Vss 0.00550397f
c73 69 Vss 0.00508271f
c74 66 Vss 0.00601821f
c75 65 Vss 3.90863e-19
c76 57 Vss 9.08254e-19
c77 56 Vss 6.01198e-19
c78 54 Vss 0.00400006f
c79 51 Vss 0.00786937f
c80 49 Vss 0.135055f
c81 45 Vss 0.127825f
c82 44 Vss 9.84889e-20
c83 24 Vss 0.21954f
c84 21 Vss 0.129208f
c85 19 Vss 0.0247918f
c86 7 Vss 1.22248f
c87 4 Vss 0.139574f
r88 65 74 1.16709
r89 65 66 0.531835
r90 62 69 1.16709
r91 60 62 0.0416786
r92 57 60 0.833571
r93 56 66 10.4613
r94 53 56 0.652036
r95 53 54 8.66914
r96 52 57 0.0685365
r97 51 54 0.652036
r98 51 52 10.2113
r99 47 49 4.53833
r100 44 74 0.0238214
r101 44 45 2.26917
r102 41 44 2.26917
r103 36 49 0.00605528
r104 35 45 0.00605528
r105 32 47 0.00605528
r106 31 41 0.00605528
r107 27 69 0.0952857
r108 25 27 0.326018
r109 25 27 0.1167
r110 24 28 0.652036
r111 24 27 6.7686
r112 21 27 0.3335
r113 19 27 0.326018
r114 19 21 0.2334
r115 11 36 3.8511
r116 11 32 3.8511
r117 7 11 15.4044
r118 7 35 3.8511
r119 7 11 15.4044
r120 7 31 3.8511
r121 4 28 3.8511
r122 2 21 3.6177
.ends

.subckt PM_G5_XOR3_N2_BI 2 4 6 8 18 21 29 32 37 42 51 56 65 71 72 80 Vss
c67 80 Vss 3.59704e-19
c68 72 Vss 1.29652e-19
c69 71 Vss 7.91966e-19
c70 65 Vss 0.00113976f
c71 56 Vss 0.00255458f
c72 51 Vss 0.00236417f
c73 42 Vss 0.00116078f
c74 37 Vss 0.00223673f
c75 32 Vss 0.00202587f
c76 29 Vss 0.00450527f
c77 21 Vss 0.111942f
c78 6 Vss 0.112114f
c79 4 Vss 0.00143442f
r80 76 80 0.655813
r81 71 72 0.655813
r82 70 71 3.501
r83 65 70 0.655813
r84 42 56 1.16709
r85 42 72 2.00578
r86 37 51 1.16709
r87 37 80 12.0712
r88 37 65 2.00578
r89 32 76 2.45904
r90 29 32 1.16709
r91 21 56 0.50025
r92 18 51 0.50025
r93 8 21 3.09255
r94 6 18 3.09255
r95 4 29 0.185659
r96 2 29 0.185659
.ends

.subckt PM_G5_XOR3_N2_AI 2 4 7 11 31 37 43 46 51 60 73 79 Vss
c46 79 Vss 2.59226e-19
c47 73 Vss 0.00489127f
c48 60 Vss 0.00532163f
c49 51 Vss 0.00226804f
c50 46 Vss 0.00262268f
c51 43 Vss 0.00448639f
c52 37 Vss 0.127877f
c53 31 Vss 0.131547f
c54 7 Vss 1.20882f
c55 4 Vss 0.00143442f
r56 75 79 0.652036
r57 73 79 13.7539
r58 51 60 1.16709
r59 51 73 2.75079
r60 46 75 5.2515
r61 43 46 1.16709
r62 36 60 0.0238214
r63 36 37 2.334
r64 33 36 2.20433
r65 29 31 4.53833
r66 26 37 0.00605528
r67 25 31 0.00605528
r68 22 33 0.00605528
r69 21 29 0.00605528
r70 11 26 3.8511
r71 11 22 3.8511
r72 7 11 15.4044
r73 7 25 3.8511
r74 7 11 15.4044
r75 7 21 3.8511
r76 4 43 0.185659
r77 2 43 0.185659
.ends

.subckt PM_G5_XOR3_N2_B 2 4 6 8 16 17 24 26 33 38 42 45 50 55 60 65 73 74 80 86
+ 91 92 Vss
c75 92 Vss 1.50842e-19
c76 91 Vss 6.9543e-19
c77 86 Vss 8.71217e-19
c78 80 Vss 6.55917e-19
c79 74 Vss 5.2356e-19
c80 73 Vss 0.00528129f
c81 65 Vss 0.00250661f
c82 60 Vss 0.00217314f
c83 55 Vss 0.00427742f
c84 50 Vss 0.00149379f
c85 45 Vss 3.19996e-19
c86 42 Vss 4.98048e-19
c87 38 Vss 6.6601e-19
c88 33 Vss 1.05421e-19
c89 26 Vss 0.111942f
c90 24 Vss 9.84889e-20
c91 20 Vss 0.0247918f
c92 17 Vss 0.0339811f
c93 16 Vss 0.183683f
c94 8 Vss 0.111942f
c95 4 Vss 0.12597f
c96 2 Vss 0.136912f
r97 90 92 0.655813
r98 90 91 3.501
r99 86 91 0.655813
r100 73 80 0.0685365
r101 73 74 10.3363
r102 69 74 0.652036
r103 50 65 1.16709
r104 50 92 2.00578
r105 45 60 1.16709
r106 45 86 2.00578
r107 45 80 2.04225
r108 38 55 1.16709
r109 38 69 2.25064
r110 38 42 0.0364688
r111 36 55 0.0476429
r112 33 65 0.50025
r113 26 60 0.50025
r114 24 55 0.357321
r115 20 36 0.326018
r116 20 24 0.40845
r117 17 36 6.7686
r118 16 36 0.326018
r119 16 36 0.1167
r120 13 17 0.652036
r121 8 33 3.09255
r122 6 26 3.09255
r123 4 24 3.44265
r124 2 13 3.8511
.ends

.subckt PM_G5_XOR3_N2_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00368262f
c33 27 Vss 0.00842339f
c34 23 Vss 0.00745376f
c35 8 Vss 0.00143442f
c36 6 Vss 0.00334862f
r37 33 35 5.20982
r38 30 40 1.16709
r39 30 33 5.79332
r40 27 35 1.16709
r41 23 40 0.05
r42 8 27 0.185659
r43 6 23 0.185659
r44 4 27 0.185659
r45 2 23 0.185659
.ends

.subckt G5_XOR3_N2  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI15.X0 N_CI_XI15.X0_D N_VSS_XI15.X0_PGD N_C_XI15.X0_CG N_VSS_XI15.X0_PGD
+ N_VDD_XI15.X0_S TIGFET_HPNW8
XI12.X0 N_CI_XI12.X0_D N_VDD_XI12.X0_PGD N_C_XI12.X0_CG N_VDD_XI12.X0_PGD
+ N_VSS_XI12.X0_S TIGFET_HPNW8
XI11.X0 N_BI_XI11.X0_D N_VDD_XI11.X0_PGD N_B_XI11.X0_CG N_VDD_XI11.X0_PGD
+ N_VSS_XI11.X0_S TIGFET_HPNW8
XI13.X0 N_AI_XI13.X0_D N_VSS_XI13.X0_PGD N_A_XI13.X0_CG N_VSS_XI13.X0_PGD
+ N_VDD_XI13.X0_S TIGFET_HPNW8
XI14.X0 N_BI_XI14.X0_D N_VSS_XI14.X0_PGD N_B_XI14.X0_CG N_VSS_XI14.X0_PGD
+ N_VDD_XI14.X0_S TIGFET_HPNW8
XI0.X0 N_AI_XI0.X0_D N_VDD_XI0.X0_PGD N_A_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW8
XI18.X0 N_Z_XI18.X0_D N_AI_XI18.X0_PGD N_BI_XI18.X0_CG N_AI_XI18.X0_PGD
+ N_C_XI18.X0_S TIGFET_HPNW8
XI16.X0 N_Z_XI16.X0_D N_AI_XI16.X0_PGD N_B_XI16.X0_CG N_AI_XI16.X0_PGD
+ N_CI_XI16.X0_S TIGFET_HPNW8
XI19.X0 N_Z_XI19.X0_D N_A_XI19.X0_PGD N_B_XI19.X0_CG N_A_XI19.X0_PGD
+ N_C_XI19.X0_S TIGFET_HPNW8
XI17.X0 N_Z_XI17.X0_D N_A_XI17.X0_PGD N_BI_XI17.X0_CG N_A_XI17.X0_PGD
+ N_CI_XI17.X0_S TIGFET_HPNW8
*
x_PM_G5_XOR3_N2_VDD N_VDD_XI15.X0_S N_VDD_XI12.X0_PGD N_VDD_XI11.X0_PGD
+ N_VDD_XI13.X0_S N_VDD_XI14.X0_S N_VDD_XI0.X0_PGD N_VDD_c_112_p N_VDD_c_20_p
+ N_VDD_c_25_p N_VDD_c_4_p N_VDD_c_93_p N_VDD_c_102_p N_VDD_c_21_p N_VDD_c_75_p
+ N_VDD_c_103_p N_VDD_c_6_p N_VDD_c_7_p N_VDD_c_13_p N_VDD_c_5_p N_VDD_c_62_p
+ N_VDD_c_30_p N_VDD_c_63_p N_VDD_c_31_p N_VDD_c_17_p N_VDD_c_64_p N_VDD_c_22_p
+ N_VDD_c_10_p N_VDD_c_26_p N_VDD_c_38_p N_VDD_c_11_p N_VDD_c_58_p VDD
+ N_VDD_c_66_p N_VDD_c_70_p N_VDD_c_2_p N_VDD_c_43_p N_VDD_c_39_p Vss
+ PM_G5_XOR3_N2_VDD
x_PM_G5_XOR3_N2_C N_C_XI15.X0_CG N_C_XI12.X0_CG N_C_XI18.X0_S N_C_XI19.X0_S
+ N_C_c_134_p N_C_c_118_n N_C_c_128_p N_C_c_121_n N_C_c_165_p C N_C_c_130_p
+ N_C_c_148_p N_C_c_167_p N_C_c_124_n N_C_c_125_n N_C_c_150_p N_C_c_154_p Vss
+ PM_G5_XOR3_N2_C
x_PM_G5_XOR3_N2_VSS N_VSS_XI15.X0_PGD N_VSS_XI12.X0_S N_VSS_XI11.X0_S
+ N_VSS_XI13.X0_PGD N_VSS_XI14.X0_PGD N_VSS_XI0.X0_S N_VSS_c_179_n N_VSS_c_235_n
+ N_VSS_c_180_n N_VSS_c_182_n N_VSS_c_183_n N_VSS_c_184_n N_VSS_c_289_p
+ N_VSS_c_186_n N_VSS_c_252_p N_VSS_c_187_n N_VSS_c_192_n N_VSS_c_195_n
+ N_VSS_c_199_n N_VSS_c_203_n N_VSS_c_204_n N_VSS_c_207_n N_VSS_c_211_n
+ N_VSS_c_215_n N_VSS_c_218_n N_VSS_c_220_n N_VSS_c_221_n N_VSS_c_222_n
+ N_VSS_c_226_n N_VSS_c_227_n N_VSS_c_230_n N_VSS_c_286_p N_VSS_c_231_n
+ N_VSS_c_232_n N_VSS_c_233_n VSS Vss PM_G5_XOR3_N2_VSS
x_PM_G5_XOR3_N2_CI N_CI_XI15.X0_D N_CI_XI12.X0_D N_CI_XI16.X0_S N_CI_XI17.X0_S
+ N_CI_c_296_n N_CI_c_309_n N_CI_c_343_p N_CI_c_298_n N_CI_c_316_n N_CI_c_345_p
+ N_CI_c_302_n N_CI_c_319_n N_CI_c_320_n N_CI_c_333_p N_CI_c_326_p Vss
+ PM_G5_XOR3_N2_CI
x_PM_G5_XOR3_N2_A N_A_XI13.X0_CG N_A_XI0.X0_CG N_A_XI19.X0_PGD N_A_XI17.X0_PGD
+ N_A_c_351_n N_A_c_405_p N_A_c_396_p N_A_c_398_p N_A_c_352_n N_A_c_358_n
+ N_A_c_359_n N_A_c_360_n A N_A_c_367_n N_A_c_368_n N_A_c_361_n N_A_c_410_p Vss
+ PM_G5_XOR3_N2_A
x_PM_G5_XOR3_N2_BI N_BI_XI11.X0_D N_BI_XI14.X0_D N_BI_XI18.X0_CG N_BI_XI17.X0_CG
+ N_BI_c_446_n N_BI_c_447_n N_BI_c_423_n N_BI_c_426_n N_BI_c_430_n N_BI_c_443_n
+ N_BI_c_453_n N_BI_c_455_n N_BI_c_433_n N_BI_c_476_p N_BI_c_444_n N_BI_c_434_n
+ Vss PM_G5_XOR3_N2_BI
x_PM_G5_XOR3_N2_AI N_AI_XI13.X0_D N_AI_XI0.X0_D N_AI_XI18.X0_PGD
+ N_AI_XI16.X0_PGD N_AI_c_500_n N_AI_c_491_n N_AI_c_492_n N_AI_c_494_n
+ N_AI_c_507_n N_AI_c_530_p N_AI_c_498_n N_AI_c_510_n Vss PM_G5_XOR3_N2_AI
x_PM_G5_XOR3_N2_B N_B_XI11.X0_CG N_B_XI14.X0_CG N_B_XI16.X0_CG N_B_XI19.X0_CG
+ N_B_c_537_n N_B_c_538_n N_B_c_546_n N_B_c_600_n N_B_c_564_n N_B_c_539_n B
+ N_B_c_580_n N_B_c_554_n N_B_c_540_n N_B_c_585_n N_B_c_572_n N_B_c_541_n
+ N_B_c_556_n N_B_c_557_n N_B_c_543_n N_B_c_597_n N_B_c_544_n Vss
+ PM_G5_XOR3_N2_B
x_PM_G5_XOR3_N2_Z N_Z_XI18.X0_D N_Z_XI16.X0_D N_Z_XI19.X0_D N_Z_XI17.X0_D
+ N_Z_c_611_n N_Z_c_618_n N_Z_c_615_n Z Vss PM_G5_XOR3_N2_Z
cc_1 N_VDD_XI11.X0_PGD N_C_XI12.X0_CG 0.00111653f
cc_2 N_VDD_c_2_p N_C_XI12.X0_CG 9.52277e-19
cc_3 N_VDD_XI12.X0_PGD N_C_c_118_n 4.18724e-19
cc_4 N_VDD_c_4_p N_C_c_118_n 0.00111653f
cc_5 N_VDD_c_5_p N_C_c_118_n 0.00134893f
cc_6 N_VDD_c_6_p N_C_c_121_n 3.43419e-19
cc_7 N_VDD_c_7_p C 4.76491e-19
cc_8 N_VDD_c_5_p C 0.00161703f
cc_9 N_VDD_c_5_p N_C_c_124_n 2.84956e-19
cc_10 N_VDD_c_10_p N_C_c_125_n 4.83409e-19
cc_11 N_VDD_c_11_p N_C_c_125_n 7.93016e-19
cc_12 N_VDD_XI12.X0_PGD N_VSS_XI15.X0_PGD 0.00201307f
cc_13 N_VDD_c_13_p N_VSS_XI15.X0_PGD 3.1461e-19
cc_14 N_VDD_c_5_p N_VSS_XI15.X0_PGD 2.01827e-19
cc_15 N_VDD_XI11.X0_PGD N_VSS_XI13.X0_PGD 2.35243e-19
cc_16 N_VDD_XI0.X0_PGD N_VSS_XI13.X0_PGD 0.00201252f
cc_17 N_VDD_c_17_p N_VSS_XI13.X0_PGD 3.00522e-19
cc_18 N_VDD_XI11.X0_PGD N_VSS_XI14.X0_PGD 0.00200584f
cc_19 N_VDD_XI0.X0_PGD N_VSS_XI14.X0_PGD 2.22638e-19
cc_20 N_VDD_c_20_p N_VSS_c_179_n 0.00201307f
cc_21 N_VDD_c_21_p N_VSS_c_180_n 0.00201252f
cc_22 N_VDD_c_22_p N_VSS_c_180_n 2.84671e-19
cc_23 N_VDD_c_22_p N_VSS_c_182_n 3.9313e-19
cc_24 N_VDD_c_11_p N_VSS_c_183_n 2.41035e-19
cc_25 N_VDD_c_25_p N_VSS_c_184_n 0.00200584f
cc_26 N_VDD_c_26_p N_VSS_c_184_n 3.9313e-19
cc_27 N_VDD_c_5_p N_VSS_c_186_n 3.4118e-19
cc_28 N_VDD_c_13_p N_VSS_c_187_n 4.32468e-19
cc_29 N_VDD_c_5_p N_VSS_c_187_n 3.85027e-19
cc_30 N_VDD_c_30_p N_VSS_c_187_n 0.00120518f
cc_31 N_VDD_c_31_p N_VSS_c_187_n 3.98949e-19
cc_32 N_VDD_c_2_p N_VSS_c_187_n 3.48267e-19
cc_33 N_VDD_c_5_p N_VSS_c_192_n 3.98099e-19
cc_34 N_VDD_c_10_p N_VSS_c_192_n 7.43603e-19
cc_35 N_VDD_c_11_p N_VSS_c_192_n 5.11768e-19
cc_36 N_VDD_c_17_p N_VSS_c_195_n 6.74818e-19
cc_37 N_VDD_c_22_p N_VSS_c_195_n 0.00161703f
cc_38 N_VDD_c_38_p N_VSS_c_195_n 8.6926e-19
cc_39 N_VDD_c_39_p N_VSS_c_195_n 3.48267e-19
cc_40 N_VDD_c_10_p N_VSS_c_199_n 6.78479e-19
cc_41 N_VDD_c_26_p N_VSS_c_199_n 0.00161703f
cc_42 N_VDD_c_11_p N_VSS_c_199_n 0.00242479f
cc_43 N_VDD_c_43_p N_VSS_c_199_n 3.48267e-19
cc_44 N_VDD_c_38_p N_VSS_c_203_n 7.32365e-19
cc_45 N_VDD_c_13_p N_VSS_c_204_n 4.41003e-19
cc_46 N_VDD_c_31_p N_VSS_c_204_n 3.89161e-19
cc_47 N_VDD_c_2_p N_VSS_c_204_n 7.99831e-19
cc_48 N_VDD_c_17_p N_VSS_c_207_n 3.48267e-19
cc_49 N_VDD_c_22_p N_VSS_c_207_n 2.26455e-19
cc_50 N_VDD_c_38_p N_VSS_c_207_n 3.99794e-19
cc_51 N_VDD_c_39_p N_VSS_c_207_n 6.489e-19
cc_52 N_VDD_c_10_p N_VSS_c_211_n 3.82294e-19
cc_53 N_VDD_c_26_p N_VSS_c_211_n 2.26455e-19
cc_54 N_VDD_c_11_p N_VSS_c_211_n 9.55109e-19
cc_55 N_VDD_c_43_p N_VSS_c_211_n 6.46219e-19
cc_56 N_VDD_c_7_p N_VSS_c_215_n 0.00347459f
cc_57 N_VDD_c_13_p N_VSS_c_215_n 0.00229697f
cc_58 N_VDD_c_58_p N_VSS_c_215_n 0.0010705f
cc_59 N_VDD_c_13_p N_VSS_c_218_n 0.0086177f
cc_60 N_VDD_c_31_p N_VSS_c_218_n 0.00116809f
cc_61 N_VDD_c_5_p N_VSS_c_220_n 0.00954271f
cc_62 N_VDD_c_62_p N_VSS_c_221_n 0.00107367f
cc_63 N_VDD_c_63_p N_VSS_c_222_n 0.00827847f
cc_64 N_VDD_c_64_p N_VSS_c_222_n 7.30484e-19
cc_65 N_VDD_c_22_p N_VSS_c_222_n 0.00369102f
cc_66 N_VDD_c_66_p N_VSS_c_222_n 0.00149929f
cc_67 N_VDD_c_13_p N_VSS_c_226_n 0.0010758f
cc_68 N_VDD_c_5_p N_VSS_c_227_n 0.00143208f
cc_69 N_VDD_c_26_p N_VSS_c_227_n 0.00601868f
cc_70 N_VDD_c_70_p N_VSS_c_227_n 0.00107091f
cc_71 N_VDD_c_22_p N_VSS_c_230_n 0.00534674f
cc_72 N_VDD_c_13_p N_VSS_c_231_n 0.00112682f
cc_73 N_VDD_c_5_p N_VSS_c_232_n 0.00107375f
cc_74 N_VDD_c_22_p N_VSS_c_233_n 7.74609e-19
cc_75 N_VDD_c_75_p N_CI_c_296_n 3.43419e-19
cc_76 N_VDD_c_30_p N_CI_c_296_n 3.72199e-19
cc_77 N_VDD_c_75_p N_CI_c_298_n 3.48267e-19
cc_78 N_VDD_c_5_p N_CI_c_298_n 4.34701e-19
cc_79 N_VDD_c_30_p N_CI_c_298_n 5.226e-19
cc_80 N_VDD_c_31_p N_CI_c_298_n 0.00101464f
cc_81 N_VDD_c_31_p N_CI_c_302_n 6.82638e-19
cc_82 N_VDD_c_64_p N_CI_c_302_n 7.0762e-19
cc_83 N_VDD_XI0.X0_PGD N_A_c_351_n 3.94784e-19
cc_84 N_VDD_XI0.X0_PGD N_A_c_352_n 2.73656e-19
cc_85 N_VDD_c_6_p N_A_c_352_n 2.69869e-19
cc_86 N_VDD_c_22_p N_A_c_352_n 4.57714e-19
cc_87 N_VDD_c_38_p N_A_c_352_n 3.99109e-19
cc_88 N_VDD_c_11_p N_A_c_352_n 3.90005e-19
cc_89 N_VDD_c_39_p N_A_c_352_n 2.43883e-19
cc_90 N_VDD_c_6_p N_A_c_358_n 9.18655e-19
cc_91 N_VDD_c_11_p N_A_c_359_n 0.00564482f
cc_92 N_VDD_c_31_p N_A_c_360_n 0.00104501f
cc_93 N_VDD_c_93_p N_A_c_361_n 3.61944e-19
cc_94 N_VDD_c_31_p N_A_c_361_n 5.71421e-19
cc_95 N_VDD_c_6_p N_BI_c_423_n 3.43419e-19
cc_96 N_VDD_c_26_p N_BI_c_423_n 3.4118e-19
cc_97 N_VDD_c_11_p N_BI_c_423_n 3.48267e-19
cc_98 N_VDD_c_6_p N_BI_c_426_n 3.48267e-19
cc_99 N_VDD_c_26_p N_BI_c_426_n 3.98099e-19
cc_100 N_VDD_c_11_p N_BI_c_426_n 4.99861e-19
cc_101 N_VDD_XI0.X0_PGD N_AI_XI18.X0_PGD 3.2392e-19
cc_102 N_VDD_c_102_p N_AI_c_491_n 3.2392e-19
cc_103 N_VDD_c_103_p N_AI_c_492_n 3.43419e-19
cc_104 N_VDD_c_64_p N_AI_c_492_n 3.73302e-19
cc_105 N_VDD_c_103_p N_AI_c_494_n 3.48267e-19
cc_106 N_VDD_c_64_p N_AI_c_494_n 5.23123e-19
cc_107 N_VDD_c_22_p N_AI_c_494_n 4.34701e-19
cc_108 N_VDD_c_38_p N_AI_c_494_n 5.44192e-19
cc_109 N_VDD_c_22_p N_AI_c_498_n 4.11874e-19
cc_110 N_VDD_XI12.X0_PGD N_B_XI11.X0_CG 0.00111821f
cc_111 N_VDD_XI11.X0_PGD N_B_c_537_n 3.99339e-19
cc_112 N_VDD_c_112_p N_B_c_538_n 0.00111821f
cc_113 N_VDD_c_31_p N_B_c_539_n 7.52847e-19
cc_114 N_VDD_c_39_p N_B_c_540_n 4.92948e-19
cc_115 N_VDD_c_11_p N_B_c_541_n 3.15013e-19
cc_116 N_C_c_118_n N_VSS_XI15.X0_PGD 4.18724e-19
cc_117 N_C_c_128_p N_VSS_c_235_n 4.96533e-19
cc_118 C N_VSS_c_187_n 2.70019e-19
cc_119 N_C_c_130_p N_VSS_c_187_n 2.56587e-19
cc_120 N_C_c_125_n N_VSS_c_187_n 2.07529e-19
cc_121 N_C_c_125_n N_VSS_c_192_n 0.00194391f
cc_122 N_C_c_125_n N_VSS_c_199_n 0.00158941f
cc_123 N_C_c_134_p N_VSS_c_204_n 0.00249737f
cc_124 C N_VSS_c_204_n 2.87758e-19
cc_125 N_C_c_124_n N_VSS_c_204_n 2.0363e-19
cc_126 N_C_c_130_p N_VSS_c_215_n 4.01014e-19
cc_127 N_C_c_125_n N_VSS_c_215_n 2.67374e-19
cc_128 C N_VSS_c_220_n 3.52403e-19
cc_129 N_C_c_130_p N_VSS_c_220_n 0.00136475f
cc_130 N_C_c_125_n N_VSS_c_220_n 0.00317947f
cc_131 N_C_c_125_n N_VSS_c_227_n 0.00191592f
cc_132 N_C_c_118_n N_CI_c_296_n 6.55689e-19
cc_133 N_C_c_125_n N_CI_c_298_n 0.00101026f
cc_134 N_C_c_125_n N_CI_c_302_n 0.00289054f
cc_135 N_C_c_125_n N_A_c_352_n 2.24413e-19
cc_136 N_C_c_121_n N_A_c_358_n 8.20481e-19
cc_137 N_C_c_148_p N_A_c_358_n 0.00195474f
cc_138 N_C_c_125_n N_A_c_359_n 4.776e-19
cc_139 N_C_c_150_p N_A_c_367_n 2.7748e-19
cc_140 N_C_c_148_p N_A_c_368_n 0.0018313f
cc_141 N_C_c_125_n N_A_c_368_n 3.28319e-19
cc_142 N_C_c_150_p N_A_c_368_n 0.00220096f
cc_143 N_C_c_154_p N_A_c_368_n 2.81326e-19
cc_144 N_C_c_125_n N_BI_c_426_n 0.00113193f
cc_145 N_C_c_148_p N_BI_c_430_n 0.00119554f
cc_146 N_C_c_125_n N_BI_c_430_n 0.00400118f
cc_147 N_C_c_150_p N_BI_c_430_n 6.70289e-19
cc_148 N_C_c_150_p N_BI_c_433_n 8.45766e-19
cc_149 N_C_c_125_n N_BI_c_434_n 6.63379e-19
cc_150 N_C_c_148_p N_B_c_541_n 4.44753e-19
cc_151 N_C_c_150_p N_B_c_543_n 3.99616e-19
cc_152 N_C_c_150_p N_B_c_544_n 0.00180761f
cc_153 N_C_c_121_n N_Z_c_611_n 3.43419e-19
cc_154 N_C_c_165_p N_Z_c_611_n 3.43419e-19
cc_155 N_C_c_148_p N_Z_c_611_n 3.48267e-19
cc_156 N_C_c_167_p N_Z_c_611_n 3.48267e-19
cc_157 N_C_c_165_p N_Z_c_615_n 3.48267e-19
cc_158 N_C_c_148_p N_Z_c_615_n 6.09821e-19
cc_159 N_C_c_167_p N_Z_c_615_n 5.71987e-19
cc_160 N_VSS_c_186_n N_CI_c_296_n 3.43419e-19
cc_161 N_VSS_c_192_n N_CI_c_296_n 3.48267e-19
cc_162 N_VSS_c_252_p N_CI_c_309_n 3.43419e-19
cc_163 N_VSS_c_186_n N_CI_c_298_n 3.48267e-19
cc_164 N_VSS_c_187_n N_CI_c_298_n 5.88914e-19
cc_165 N_VSS_c_192_n N_CI_c_298_n 8.10527e-19
cc_166 N_VSS_c_215_n N_CI_c_298_n 4.71364e-19
cc_167 N_VSS_c_218_n N_CI_c_298_n 9.66309e-19
cc_168 N_VSS_c_220_n N_CI_c_298_n 2.82247e-19
cc_169 N_VSS_c_203_n N_CI_c_316_n 8.74405e-19
cc_170 N_VSS_c_195_n N_CI_c_302_n 3.79792e-19
cc_171 N_VSS_c_230_n N_CI_c_302_n 5.41979e-19
cc_172 N_VSS_c_222_n N_CI_c_319_n 0.00182487f
cc_173 N_VSS_c_203_n N_CI_c_320_n 0.00142004f
cc_174 N_VSS_XI13.X0_PGD N_A_c_351_n 3.91587e-19
cc_175 N_VSS_c_203_n N_A_c_352_n 8.4508e-19
cc_176 N_VSS_c_230_n N_A_c_352_n 4.69076e-19
cc_177 N_VSS_c_195_n N_A_c_360_n 3.32273e-19
cc_178 N_VSS_c_207_n N_A_c_360_n 3.1261e-19
cc_179 N_VSS_c_195_n N_A_c_361_n 3.04912e-19
cc_180 N_VSS_c_207_n N_A_c_361_n 0.00110478f
cc_181 N_VSS_c_186_n N_BI_c_423_n 3.43419e-19
cc_182 N_VSS_c_192_n N_BI_c_423_n 3.48267e-19
cc_183 N_VSS_c_186_n N_BI_c_426_n 3.48267e-19
cc_184 N_VSS_c_192_n N_BI_c_426_n 8.10527e-19
cc_185 N_VSS_c_227_n N_BI_c_426_n 2.79692e-19
cc_186 N_VSS_XI14.X0_PGD N_AI_XI18.X0_PGD 2.74627e-19
cc_187 N_VSS_c_183_n N_AI_c_500_n 2.74627e-19
cc_188 N_VSS_c_252_p N_AI_c_492_n 3.43419e-19
cc_189 N_VSS_c_203_n N_AI_c_492_n 3.48267e-19
cc_190 N_VSS_c_252_p N_AI_c_494_n 3.48267e-19
cc_191 N_VSS_c_195_n N_AI_c_494_n 0.00108072f
cc_192 N_VSS_c_203_n N_AI_c_494_n 0.00213737f
cc_193 N_VSS_c_230_n N_AI_c_494_n 2.86662e-19
cc_194 N_VSS_c_203_n N_AI_c_507_n 0.00122373f
cc_195 N_VSS_c_230_n N_AI_c_498_n 0.00370204f
cc_196 N_VSS_c_286_p N_AI_c_498_n 0.0017148f
cc_197 N_VSS_c_230_n N_AI_c_510_n 0.0018958f
cc_198 N_VSS_XI14.X0_PGD N_B_c_537_n 3.96142e-19
cc_199 N_VSS_c_289_p N_B_c_546_n 9.56171e-19
cc_200 N_VSS_c_199_n N_B_c_539_n 2.57202e-19
cc_201 N_VSS_c_199_n B 3.42746e-19
cc_202 N_VSS_c_211_n B 3.2351e-19
cc_203 N_VSS_c_199_n N_B_c_540_n 3.2351e-19
cc_204 N_VSS_c_211_n N_B_c_540_n 2.68747e-19
cc_205 N_VSS_c_203_n N_B_c_541_n 3.58501e-19
cc_206 N_CI_c_302_n N_A_c_352_n 0.00183351f
cc_207 N_CI_c_302_n N_A_c_360_n 3.36095e-19
cc_208 N_CI_c_298_n N_BI_c_426_n 9.23808e-19
cc_209 N_CI_c_316_n N_BI_c_430_n 2.81279e-19
cc_210 N_CI_c_302_n N_BI_c_430_n 0.0032559f
cc_211 N_CI_c_326_p N_BI_c_443_n 8.83269e-19
cc_212 N_CI_c_326_p N_BI_c_444_n 2.18743e-19
cc_213 N_CI_c_302_n N_BI_c_434_n 0.00153557f
cc_214 N_CI_c_302_n N_AI_c_494_n 0.00135858f
cc_215 N_CI_c_320_n N_AI_c_494_n 0.00128778f
cc_216 N_CI_c_326_p N_AI_c_507_n 0.00144463f
cc_217 N_CI_c_302_n N_AI_c_498_n 0.00198979f
cc_218 N_CI_c_333_p N_AI_c_498_n 0.00533258f
cc_219 N_CI_c_326_p N_AI_c_498_n 0.00290048f
cc_220 N_CI_c_298_n N_B_c_539_n 5.51453e-19
cc_221 N_CI_c_326_p N_B_c_554_n 6.37546e-19
cc_222 N_CI_c_316_n N_B_c_541_n 5.58533e-19
cc_223 N_CI_c_302_n N_B_c_556_n 0.00108926f
cc_224 N_CI_c_326_p N_B_c_557_n 2.05643e-19
cc_225 N_CI_c_302_n N_B_c_543_n 4.54861e-19
cc_226 N_CI_c_326_p N_B_c_543_n 0.00179506f
cc_227 N_CI_c_309_n N_Z_c_618_n 3.43419e-19
cc_228 N_CI_c_343_p N_Z_c_618_n 3.43419e-19
cc_229 N_CI_c_316_n N_Z_c_618_n 3.48267e-19
cc_230 N_CI_c_345_p N_Z_c_618_n 3.48267e-19
cc_231 N_CI_c_309_n N_Z_c_615_n 3.48267e-19
cc_232 N_CI_c_343_p N_Z_c_615_n 3.48267e-19
cc_233 N_CI_c_316_n N_Z_c_615_n 5.71987e-19
cc_234 N_CI_c_345_p N_Z_c_615_n 5.71987e-19
cc_235 N_CI_c_302_n N_Z_c_615_n 4.15391e-19
cc_236 N_A_c_368_n N_BI_c_446_n 2.74063e-19
cc_237 N_A_XI19.X0_PGD N_BI_c_447_n 9.65637e-19
cc_238 N_A_c_352_n N_BI_c_426_n 3.85685e-19
cc_239 N_A_c_358_n N_BI_c_426_n 4.22951e-19
cc_240 N_A_c_358_n N_BI_c_430_n 0.00110458f
cc_241 N_A_c_368_n N_BI_c_430_n 8.05288e-19
cc_242 N_A_c_368_n N_BI_c_443_n 2.98812e-19
cc_243 N_A_c_358_n N_BI_c_453_n 3.37713e-19
cc_244 N_A_c_368_n N_BI_c_453_n 2.96819e-19
cc_245 N_A_XI19.X0_PGD N_BI_c_455_n 0.00133285f
cc_246 N_A_c_368_n N_BI_c_433_n 0.00102169f
cc_247 N_A_c_352_n N_BI_c_434_n 4.10091e-19
cc_248 N_A_XI19.X0_PGD N_AI_XI18.X0_PGD 0.0174244f
cc_249 N_A_c_358_n N_AI_XI18.X0_PGD 9.55469e-19
cc_250 N_A_c_368_n N_AI_XI18.X0_PGD 7.53964e-19
cc_251 N_A_c_396_p N_AI_c_500_n 0.00199315f
cc_252 N_A_c_368_n N_AI_c_500_n 0.00125772f
cc_253 N_A_c_398_p N_AI_c_491_n 0.00201004f
cc_254 N_A_c_351_n N_AI_c_492_n 6.89066e-19
cc_255 N_A_c_352_n N_AI_c_494_n 7.80381e-19
cc_256 N_A_XI19.X0_PGD N_B_XI19.X0_CG 9.65637e-19
cc_257 N_A_c_351_n N_B_c_537_n 0.0035308f
cc_258 N_A_c_352_n N_B_c_537_n 6.06747e-19
cc_259 N_A_c_361_n N_B_c_538_n 5.83549e-19
cc_260 N_A_c_405_p N_B_c_564_n 9.37683e-19
cc_261 N_A_c_358_n N_B_c_539_n 6.35249e-19
cc_262 N_A_c_352_n B 9.05205e-19
cc_263 N_A_c_358_n B 5.05926e-19
cc_264 N_A_c_367_n N_B_c_554_n 5.53953e-19
cc_265 N_A_c_410_p N_B_c_554_n 3.2351e-19
cc_266 N_A_c_351_n N_B_c_540_n 9.10729e-19
cc_267 N_A_c_358_n N_B_c_540_n 6.84646e-19
cc_268 N_A_XI19.X0_PGD N_B_c_572_n 0.00133285f
cc_269 N_A_c_410_p N_B_c_572_n 2.68747e-19
cc_270 N_A_c_352_n N_B_c_541_n 0.00336092f
cc_271 N_A_c_358_n N_B_c_541_n 0.00192865f
cc_272 N_A_c_368_n N_B_c_541_n 8.22275e-19
cc_273 N_A_c_352_n N_B_c_556_n 5.17628e-19
cc_274 N_A_c_368_n N_Z_c_611_n 0.00107687f
cc_275 N_A_XI19.X0_PGD N_Z_c_615_n 7.94638e-19
cc_276 N_A_c_358_n N_Z_c_615_n 0.00143807f
cc_277 N_A_c_368_n N_Z_c_615_n 0.0014359f
cc_278 N_BI_XI18.X0_CG N_AI_XI18.X0_PGD 9.47088e-19
cc_279 N_BI_c_453_n N_AI_XI18.X0_PGD 0.00133285f
cc_280 N_BI_c_430_n N_AI_c_498_n 9.24953e-19
cc_281 N_BI_c_423_n N_B_c_537_n 6.89066e-19
cc_282 N_BI_c_430_n N_B_c_539_n 0.00155724f
cc_283 N_BI_c_430_n N_B_c_580_n 6.02887e-19
cc_284 N_BI_c_444_n N_B_c_580_n 3.08318e-19
cc_285 N_BI_c_443_n N_B_c_554_n 0.0017864f
cc_286 N_BI_c_455_n N_B_c_554_n 4.56568e-19
cc_287 N_BI_c_433_n N_B_c_554_n 0.00165721f
cc_288 N_BI_c_430_n N_B_c_585_n 4.56568e-19
cc_289 N_BI_c_453_n N_B_c_585_n 0.00266356f
cc_290 N_BI_c_455_n N_B_c_585_n 7.16621e-19
cc_291 N_BI_c_453_n N_B_c_572_n 6.17967e-19
cc_292 N_BI_c_455_n N_B_c_572_n 0.00243716f
cc_293 N_BI_c_430_n N_B_c_541_n 0.00391901f
cc_294 N_BI_c_430_n N_B_c_557_n 3.07174e-19
cc_295 N_BI_c_433_n N_B_c_557_n 0.00126004f
cc_296 N_BI_c_476_p N_B_c_557_n 0.00342237f
cc_297 N_BI_c_430_n N_B_c_543_n 5.09978e-19
cc_298 N_BI_c_433_n N_B_c_543_n 7.34826e-19
cc_299 N_BI_c_444_n N_B_c_543_n 8.56575e-19
cc_300 N_BI_c_476_p N_B_c_597_n 0.00210118f
cc_301 N_BI_c_430_n N_B_c_544_n 0.00142766f
cc_302 N_BI_c_433_n N_B_c_544_n 9.32988e-19
cc_303 N_BI_c_430_n N_Z_c_615_n 0.00138952f
cc_304 N_BI_c_443_n N_Z_c_615_n 0.00138952f
cc_305 N_BI_c_453_n N_Z_c_615_n 8.66889e-19
cc_306 N_BI_c_455_n N_Z_c_615_n 8.66889e-19
cc_307 N_BI_c_433_n N_Z_c_615_n 0.00103509f
cc_308 N_BI_c_476_p N_Z_c_615_n 0.00212989f
cc_309 N_BI_c_444_n N_Z_c_615_n 0.00103331f
cc_310 N_AI_XI18.X0_PGD N_B_c_600_n 9.65637e-19
cc_311 N_AI_c_507_n N_B_c_580_n 3.6769e-19
cc_312 N_AI_c_530_p N_B_c_580_n 3.2351e-19
cc_313 N_AI_XI18.X0_PGD N_B_c_585_n 0.00133285f
cc_314 N_AI_c_507_n N_B_c_585_n 3.2351e-19
cc_315 N_AI_c_530_p N_B_c_585_n 0.00117301f
cc_316 N_AI_c_507_n N_B_c_557_n 4.82497e-19
cc_317 N_AI_XI18.X0_PGD N_Z_c_615_n 4.32017e-19
cc_318 N_B_c_580_n N_Z_c_615_n 0.00157325f
cc_319 N_B_c_554_n N_Z_c_615_n 0.00138952f
cc_320 N_B_c_572_n N_Z_c_615_n 8.66889e-19
cc_321 N_B_c_557_n N_Z_c_615_n 4.69528e-19
*
.ends
*
*
.subckt XOR3_HPNW8 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XOR3_N2
.ends
*
* File: G3_AND2_N3.pex.netlist
* Created: Tue Mar  1 10:56:10 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_AND2_N3_VSS 2 4 6 8 10 12 14 16 30 31 50 62 67 70 75 80 85 94 99
+ 108 109 113 114 119 125 127 132 133 134 136 Vss
c67 134 Vss 3.75522e-19
c68 133 Vss 3.62111e-19
c69 132 Vss 0.004799f
c70 127 Vss 0.00257088f
c71 125 Vss 0.00552282f
c72 119 Vss 0.00412002f
c73 114 Vss 8.41284e-19
c74 113 Vss 0.00175777f
c75 109 Vss 7.31223e-19
c76 108 Vss 0.00590165f
c77 99 Vss 0.00416928f
c78 94 Vss 0.00536429f
c79 85 Vss 7.10513e-22
c80 80 Vss 4.8997e-19
c81 75 Vss 0.00125499f
c82 70 Vss 0.00121927f
c83 67 Vss 0.0100822f
c84 62 Vss 0.00955849f
c85 58 Vss 0.0299311f
c86 57 Vss 0.0299311f
c87 51 Vss 0.0357161f
c88 50 Vss 0.0994129f
c89 42 Vss 0.107716f
c90 37 Vss 0.0688416f
c91 31 Vss 0.0350852f
c92 30 Vss 0.0646396f
c93 14 Vss 0.188821f
c94 12 Vss 0.189513f
c95 10 Vss 0.189371f
c96 8 Vss 0.190733f
c97 6 Vss 0.189919f
c98 4 Vss 0.190281f
c99 2 Vss 1.99696e-19
r100 132 136 0.326018
r101 131 132 5.50157
r102 127 131 0.655813
r103 126 134 0.494161
r104 125 136 0.326018
r105 125 126 10.1279
r106 121 134 0.128424
r107 120 133 0.494161
r108 119 134 0.494161
r109 119 120 10.378
r110 115 133 0.128424
r111 113 133 0.494161
r112 113 114 4.33457
r113 108 114 0.652036
r114 107 109 0.655813
r115 107 108 19.0471
r116 85 127 1.82344
r117 80 99 1.16709
r118 80 121 2.16729
r119 75 94 1.16709
r120 75 115 2.16729
r121 70 109 1.82344
r122 67 85 1.16709
r123 62 70 1.16709
r124 53 99 0.0476429
r125 51 53 1.45875
r126 50 54 0.652036
r127 50 53 1.45875
r128 47 51 0.652036
r129 43 58 0.494161
r130 42 44 0.652036
r131 42 43 2.9175
r132 39 58 0.128424
r133 38 57 0.494161
r134 37 58 0.494161
r135 37 38 2.8008
r136 34 57 0.128424
r137 33 94 0.0476429
r138 31 33 1.4004
r139 30 57 0.494161
r140 30 33 1.5171
r141 27 31 0.652036
r142 16 67 0.123773
r143 14 47 5.1348
r144 12 54 5.1348
r145 10 44 5.1348
r146 8 39 5.1348
r147 6 27 5.1348
r148 4 34 5.1348
r149 2 62 0.123773
.ends

.subckt PM_G3_AND2_N3_VDD 2 4 6 8 10 12 25 27 33 43 48 51 53 54 58 60 64 68 70
+ 74 76 78 79 85 94 Vss
c86 94 Vss 0.00463585f
c87 85 Vss 0.00402796f
c88 79 Vss 4.43941e-19
c89 76 Vss 4.52364e-19
c90 74 Vss 7.90245e-19
c91 70 Vss 0.00408718f
c92 68 Vss 0.00117255f
c93 64 Vss 0.00432275f
c94 60 Vss 0.00739867f
c95 58 Vss 0.00173558f
c96 55 Vss 0.00171371f
c97 54 Vss 0.0100369f
c98 53 Vss 0.00360598f
c99 51 Vss 0.00814794f
c100 48 Vss 0.00687623f
c101 43 Vss 0.00811526f
c102 33 Vss 0.0357902f
c103 32 Vss 0.102427f
c104 27 Vss 0.170038f
c105 25 Vss 0.0352365f
c106 12 Vss 0.190935f
c107 10 Vss 0.189512f
c108 8 Vss 0.00143493f
c109 2 Vss 0.221827f
r110 74 94 1.16709
r111 72 74 2.16729
r112 71 79 0.494161
r113 70 72 0.652036
r114 70 71 7.46046
r115 66 79 0.128424
r116 66 68 6.16843
r117 64 85 1.16709
r118 62 64 6.08507
r119 61 78 0.326018
r120 60 79 0.494161
r121 60 61 13.0037
r122 56 76 0.0828784
r123 56 58 1.82344
r124 54 62 0.652036
r125 54 55 10.0862
r126 53 78 0.326018
r127 52 76 0.551426
r128 52 53 5.50157
r129 51 76 0.551426
r130 50 55 0.652036
r131 50 51 15.046
r132 48 68 1.16709
r133 43 58 1.16709
r134 35 94 0.0476429
r135 33 35 1.45875
r136 32 36 0.652036
r137 32 35 1.45875
r138 29 33 0.652036
r139 27 85 0.428786
r140 25 27 5.3682
r141 22 25 0.652036
r142 12 36 5.1348
r143 10 29 5.1348
r144 8 48 0.123773
r145 6 48 0.123773
r146 4 43 0.123773
r147 2 22 6.3018
.ends

.subckt PM_G3_AND2_N3_A 1 2 9 20 23 28 33 Vss
c24 33 Vss 0.00369912f
c25 28 Vss 0.00225353f
c26 20 Vss 0.00104617f
c27 12 Vss 0.166756f
c28 1 Vss 0.171396f
r29 25 33 1.16709
r30 23 25 2.66743
r31 20 28 1.16709
r32 20 23 2.70911
r33 12 33 0.50025
r34 9 28 0.50025
r35 2 12 4.37625
r36 1 9 4.60965
.ends

.subckt PM_G3_AND2_N3_NET1 2 4 6 7 8 23 26 38 42 48 52 54 58 71 Vss
c52 71 Vss 0.00600165f
c53 60 Vss 2.11292e-19
c54 58 Vss 0.0011885f
c55 54 Vss 0.00636228f
c56 52 Vss 6.44544e-19
c57 48 Vss 8.20028e-19
c58 42 Vss 0.00560082f
c59 38 Vss 0.00901424f
c60 26 Vss 8.44333e-20
c61 23 Vss 0.229828f
c62 19 Vss 0.18045f
c63 17 Vss 0.0247918f
c64 8 Vss 0.193588f
c65 6 Vss 0.00143493f
r66 58 71 1.16709
r67 56 58 2.16729
r68 55 60 0.128424
r69 54 56 0.652036
r70 54 55 7.46046
r71 52 68 1.16709
r72 50 60 0.494161
r73 50 52 6.29346
r74 46 60 0.494161
r75 46 48 6.21011
r76 42 68 0.15
r77 38 48 1.16709
r78 26 71 0.0476429
r79 24 26 0.326018
r80 24 26 0.1167
r81 23 27 0.652036
r82 23 26 6.7686
r83 19 71 0.357321
r84 17 26 0.326018
r85 17 19 0.40845
r86 8 27 5.1348
r87 7 19 4.72635
r88 6 42 0.123773
r89 4 42 0.123773
r90 2 38 0.123773
.ends

.subckt PM_G3_AND2_N3_B 2 3 9 10 13 19 22 Vss
c26 19 Vss 2.97116e-19
c27 13 Vss 0.236449f
c28 10 Vss 0.0348969f
c29 9 Vss 0.287374f
c30 2 Vss 0.332764f
r31 19 22 0.0416786
r32 13 19 1.16709
r33 11 13 2.15895
r34 9 11 0.652036
r35 9 10 8.92755
r36 6 10 0.652036
r37 3 13 5.6016
r38 2 6 10.0362
.ends

.subckt PM_G3_AND2_N3_Z 2 4 13 16 Vss
c13 13 Vss 0.00498872f
c14 4 Vss 0.00143493f
r15 16 19 0.0416786
r16 13 19 1.16709
r17 4 13 0.123773
r18 2 13 0.123773
.ends

.subckt G3_AND2_N3  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI13.X0 N_NET1_XI13.X0_D N_VDD_XI13.X0_PGD N_A_XI13.X0_CG N_B_XI13.X0_PGS
+ N_VSS_XI13.X0_S TIGFET_HPNW12
XI15.X0 N_NET1_XI15.X0_D N_VSS_XI15.X0_PGD N_A_XI15.X0_CG N_VSS_XI15.X0_PGS
+ N_VDD_XI15.X0_S TIGFET_HPNW12
XI14.X0 N_NET1_XI14.X0_D N_VSS_XI14.X0_PGD N_B_XI14.X0_CG N_VSS_XI14.X0_PGS
+ N_VDD_XI14.X0_S TIGFET_HPNW12
XI12.X0 N_Z_XI12.X0_D N_VSS_XI12.X0_PGD N_NET1_XI12.X0_CG N_VSS_XI12.X0_PGS
+ N_VDD_XI12.X0_S TIGFET_HPNW12
XI11.X0 N_Z_XI11.X0_D N_VDD_XI11.X0_PGD N_NET1_XI11.X0_CG N_VDD_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW12
*
x_PM_G3_AND2_N3_VSS N_VSS_XI13.X0_S N_VSS_XI15.X0_PGD N_VSS_XI15.X0_PGS
+ N_VSS_XI14.X0_PGD N_VSS_XI14.X0_PGS N_VSS_XI12.X0_PGD N_VSS_XI12.X0_PGS
+ N_VSS_XI11.X0_S N_VSS_c_14_p N_VSS_c_15_p N_VSS_c_2_p N_VSS_c_3_p N_VSS_c_62_p
+ N_VSS_c_4_p N_VSS_c_8_p N_VSS_c_24_p N_VSS_c_63_p N_VSS_c_9_p N_VSS_c_26_p
+ N_VSS_c_5_p N_VSS_c_6_p N_VSS_c_18_p N_VSS_c_11_p N_VSS_c_19_p N_VSS_c_33_p
+ N_VSS_c_67_p N_VSS_c_28_p N_VSS_c_20_p N_VSS_c_34_p VSS Vss PM_G3_AND2_N3_VSS
x_PM_G3_AND2_N3_VDD N_VDD_XI13.X0_PGD N_VDD_XI15.X0_S N_VDD_XI14.X0_S
+ N_VDD_XI12.X0_S N_VDD_XI11.X0_PGD N_VDD_XI11.X0_PGS N_VDD_c_146_p
+ N_VDD_c_128_p N_VDD_c_69_n N_VDD_c_122_p N_VDD_c_123_p N_VDD_c_70_n
+ N_VDD_c_74_n N_VDD_c_79_n N_VDD_c_80_n N_VDD_c_81_n N_VDD_c_121_p N_VDD_c_88_n
+ N_VDD_c_96_n N_VDD_c_102_n N_VDD_c_105_n VDD N_VDD_c_106_n N_VDD_c_117_p
+ N_VDD_c_107_n Vss PM_G3_AND2_N3_VDD
x_PM_G3_AND2_N3_A N_A_XI13.X0_CG N_A_XI15.X0_CG N_A_c_160_n N_A_c_154_n A
+ N_A_c_163_n N_A_c_156_n Vss PM_G3_AND2_N3_A
x_PM_G3_AND2_N3_NET1 N_NET1_XI13.X0_D N_NET1_XI15.X0_D N_NET1_XI14.X0_D
+ N_NET1_XI12.X0_CG N_NET1_XI11.X0_CG N_NET1_c_178_n N_NET1_c_179_n
+ N_NET1_c_180_n N_NET1_c_194_n N_NET1_c_182_n N_NET1_c_185_n N_NET1_c_186_n
+ N_NET1_c_188_n N_NET1_c_190_n Vss PM_G3_AND2_N3_NET1
x_PM_G3_AND2_N3_B N_B_XI13.X0_PGS N_B_XI14.X0_CG N_B_c_230_n N_B_c_232_n
+ N_B_c_237_n N_B_c_252_n B Vss PM_G3_AND2_N3_B
x_PM_G3_AND2_N3_Z N_Z_XI12.X0_D N_Z_XI11.X0_D N_Z_c_256_n Z Vss PM_G3_AND2_N3_Z
cc_1 N_VSS_XI12.X0_PGD N_VDD_XI11.X0_PGD 0.00195824f
cc_2 N_VSS_c_2_p N_VDD_c_69_n 0.00195824f
cc_3 N_VSS_c_3_p N_VDD_c_70_n 9.5668e-19
cc_4 N_VSS_c_4_p N_VDD_c_70_n 0.00165395f
cc_5 N_VSS_c_5_p N_VDD_c_70_n 0.00795264f
cc_6 N_VSS_c_6_p N_VDD_c_70_n 0.00190019f
cc_7 N_VSS_XI15.X0_PGS N_VDD_c_74_n 3.39564e-19
cc_8 N_VSS_c_8_p N_VDD_c_74_n 4.42007e-19
cc_9 N_VSS_c_9_p N_VDD_c_74_n 3.70842e-19
cc_10 N_VSS_c_5_p N_VDD_c_74_n 0.00357958f
cc_11 N_VSS_c_11_p N_VDD_c_74_n 0.00107567f
cc_12 N_VSS_c_4_p N_VDD_c_79_n 0.00237483f
cc_13 N_VSS_c_4_p N_VDD_c_80_n 3.67743e-19
cc_14 N_VSS_c_14_p N_VDD_c_81_n 0.00161328f
cc_15 N_VSS_c_15_p N_VDD_c_81_n 3.76573e-19
cc_16 N_VSS_c_8_p N_VDD_c_81_n 0.00161703f
cc_17 N_VSS_c_9_p N_VDD_c_81_n 2.26455e-19
cc_18 N_VSS_c_18_p N_VDD_c_81_n 0.00349492f
cc_19 N_VSS_c_19_p N_VDD_c_81_n 0.00593063f
cc_20 N_VSS_c_20_p N_VDD_c_81_n 7.61747e-19
cc_21 N_VSS_XI14.X0_PGS N_VDD_c_88_n 2.0368e-19
cc_22 N_VSS_XI12.X0_PGS N_VDD_c_88_n 2.24983e-19
cc_23 N_VSS_c_8_p N_VDD_c_88_n 6.58919e-19
cc_24 N_VSS_c_24_p N_VDD_c_88_n 0.0018079f
cc_25 N_VSS_c_9_p N_VDD_c_88_n 2.56577e-19
cc_26 N_VSS_c_26_p N_VDD_c_88_n 9.55109e-19
cc_27 N_VSS_c_5_p N_VDD_c_88_n 4.30333e-19
cc_28 N_VSS_c_28_p N_VDD_c_88_n 2.91233e-19
cc_29 N_VSS_c_2_p N_VDD_c_96_n 5.15102e-19
cc_30 N_VSS_c_24_p N_VDD_c_96_n 0.00161703f
cc_31 N_VSS_c_26_p N_VDD_c_96_n 2.26455e-19
cc_32 N_VSS_c_19_p N_VDD_c_96_n 0.00133474f
cc_33 N_VSS_c_33_p N_VDD_c_96_n 0.00600556f
cc_34 N_VSS_c_34_p N_VDD_c_96_n 7.74609e-19
cc_35 N_VSS_c_24_p N_VDD_c_102_n 8.50587e-19
cc_36 N_VSS_c_26_p N_VDD_c_102_n 3.82294e-19
cc_37 N_VSS_c_28_p N_VDD_c_102_n 3.85245e-19
cc_38 N_VSS_c_5_p N_VDD_c_105_n 0.00100712f
cc_39 N_VSS_c_19_p N_VDD_c_106_n 9.82771e-19
cc_40 N_VSS_c_24_p N_VDD_c_107_n 3.48267e-19
cc_41 N_VSS_c_26_p N_VDD_c_107_n 6.46219e-19
cc_42 N_VSS_c_9_p N_A_c_154_n 2.354e-19
cc_43 N_VSS_c_5_p N_A_c_154_n 0.00149458f
cc_44 N_VSS_c_8_p N_A_c_156_n 2.15082e-19
cc_45 N_VSS_c_9_p N_A_c_156_n 4.9359e-19
cc_46 N_VSS_XI12.X0_PGD N_NET1_c_178_n 4.31283e-19
cc_47 N_VSS_c_26_p N_NET1_c_179_n 5.28949e-19
cc_48 N_VSS_c_3_p N_NET1_c_180_n 3.43419e-19
cc_49 N_VSS_c_4_p N_NET1_c_180_n 3.48267e-19
cc_50 N_VSS_c_3_p N_NET1_c_182_n 3.48267e-19
cc_51 N_VSS_c_4_p N_NET1_c_182_n 8.50248e-19
cc_52 N_VSS_c_5_p N_NET1_c_182_n 8.95101e-19
cc_53 N_VSS_c_19_p N_NET1_c_185_n 2.278e-19
cc_54 N_VSS_XI14.X0_PGS N_NET1_c_186_n 2.25423e-19
cc_55 N_VSS_c_19_p N_NET1_c_186_n 4.57847e-19
cc_56 N_VSS_c_24_p N_NET1_c_188_n 2.00623e-19
cc_57 N_VSS_c_26_p N_NET1_c_188_n 2.28697e-19
cc_58 N_VSS_c_24_p N_NET1_c_190_n 2.15082e-19
cc_59 N_VSS_XI15.X0_PGD N_B_c_230_n 8.16475e-19
cc_60 N_VSS_XI14.X0_PGD N_B_c_230_n 8.16475e-19
cc_61 N_VSS_XI15.X0_PGS N_B_c_232_n 0.00101175f
cc_62 N_VSS_c_62_p N_Z_c_256_n 3.43419e-19
cc_63 N_VSS_c_63_p N_Z_c_256_n 3.48267e-19
cc_64 N_VSS_c_62_p Z 3.48267e-19
cc_65 N_VSS_c_63_p Z 4.99861e-19
cc_66 N_VSS_c_33_p Z 2.23989e-19
cc_67 N_VSS_c_67_p Z 2.7826e-19
cc_68 N_VDD_XI13.X0_PGD N_A_XI13.X0_CG 4.85665e-19
cc_69 N_VDD_c_79_n N_A_XI13.X0_CG 3.10124e-19
cc_70 N_VDD_c_79_n N_A_c_160_n 2.67445e-19
cc_71 N_VDD_c_70_n N_A_c_154_n 0.0028804f
cc_72 N_VDD_c_79_n N_A_c_154_n 4.70376e-19
cc_73 N_VDD_XI13.X0_PGD N_A_c_163_n 4.86892e-19
cc_74 N_VDD_c_70_n N_A_c_163_n 3.66936e-19
cc_75 N_VDD_c_79_n N_A_c_163_n 2.64879e-19
cc_76 N_VDD_c_117_p N_A_c_163_n 5.21476e-19
cc_77 N_VDD_c_70_n N_A_c_156_n 5.07754e-19
cc_78 N_VDD_XI11.X0_PGD N_NET1_c_178_n 4.31283e-19
cc_79 N_VDD_c_79_n N_NET1_c_180_n 0.0011619f
cc_80 N_VDD_c_121_p N_NET1_c_180_n 8.835e-19
cc_81 N_VDD_c_122_p N_NET1_c_194_n 3.43419e-19
cc_82 N_VDD_c_123_p N_NET1_c_194_n 3.43419e-19
cc_83 N_VDD_c_80_n N_NET1_c_194_n 3.72199e-19
cc_84 N_VDD_c_81_n N_NET1_c_194_n 2.82909e-19
cc_85 N_VDD_c_88_n N_NET1_c_194_n 3.48267e-19
cc_86 N_VDD_XI13.X0_PGD N_NET1_c_182_n 3.17068e-19
cc_87 N_VDD_c_128_p N_NET1_c_182_n 8.01918e-19
cc_88 N_VDD_c_70_n N_NET1_c_182_n 0.00133415f
cc_89 N_VDD_c_79_n N_NET1_c_182_n 0.00168724f
cc_90 N_VDD_c_121_p N_NET1_c_182_n 0.00619213f
cc_91 N_VDD_c_117_p N_NET1_c_182_n 9.07013e-19
cc_92 N_VDD_c_122_p N_NET1_c_185_n 3.48267e-19
cc_93 N_VDD_c_123_p N_NET1_c_185_n 3.48267e-19
cc_94 N_VDD_c_80_n N_NET1_c_185_n 8.08807e-19
cc_95 N_VDD_c_81_n N_NET1_c_185_n 3.96039e-19
cc_96 N_VDD_c_88_n N_NET1_c_185_n 7.82265e-19
cc_97 N_VDD_c_128_p N_NET1_c_186_n 3.89384e-19
cc_98 N_VDD_c_123_p N_NET1_c_186_n 2.74986e-19
cc_99 N_VDD_c_121_p N_NET1_c_186_n 0.00138769f
cc_100 N_VDD_c_88_n N_NET1_c_186_n 5.47694e-19
cc_101 N_VDD_c_117_p N_NET1_c_186_n 8.66889e-19
cc_102 N_VDD_XI13.X0_PGD N_B_XI13.X0_PGS 0.00331493f
cc_103 N_VDD_c_70_n N_B_XI13.X0_PGS 7.63549e-19
cc_104 N_VDD_c_79_n N_B_XI13.X0_PGS 6.44483e-19
cc_105 N_VDD_c_146_p N_B_c_230_n 0.00792574f
cc_106 N_VDD_c_117_p N_B_c_237_n 0.0014275f
cc_107 N_VDD_c_123_p N_Z_c_256_n 3.43419e-19
cc_108 N_VDD_c_88_n N_Z_c_256_n 3.48267e-19
cc_109 N_VDD_c_96_n N_Z_c_256_n 2.74986e-19
cc_110 N_VDD_c_123_p Z 3.48267e-19
cc_111 N_VDD_c_88_n Z 7.09569e-19
cc_112 N_VDD_c_96_n Z 3.66281e-19
cc_113 N_A_c_154_n N_NET1_c_182_n 0.0080879f
cc_114 N_A_c_163_n N_NET1_c_182_n 8.85473e-19
cc_115 N_A_c_156_n N_NET1_c_185_n 9.58642e-19
cc_116 N_A_XI13.X0_CG N_B_XI13.X0_PGS 4.84447e-19
cc_117 N_A_c_154_n N_B_XI13.X0_PGS 3.59952e-19
cc_118 N_A_c_163_n N_B_XI13.X0_PGS 5.64689e-19
cc_119 N_A_c_154_n N_B_c_230_n 2.067e-19
cc_120 N_A_c_163_n N_B_c_230_n 6.90429e-19
cc_121 N_A_c_156_n N_B_c_230_n 0.0015879f
cc_122 N_A_c_156_n N_B_c_237_n 9.27569e-19
cc_123 N_NET1_c_194_n N_B_c_230_n 3.4562e-19
cc_124 N_NET1_c_185_n N_B_c_230_n 2.39796e-19
cc_125 N_NET1_c_186_n N_B_c_230_n 4.12724e-19
cc_126 N_NET1_c_185_n N_B_c_237_n 0.00116203f
cc_127 N_NET1_c_186_n N_B_c_237_n 0.00112058f
cc_128 N_NET1_c_188_n N_B_c_237_n 3.86148e-19
cc_129 N_NET1_c_190_n N_B_c_237_n 0.00196155f
cc_130 N_NET1_c_185_n N_B_c_252_n 0.00147455f
cc_131 N_NET1_c_186_n N_B_c_252_n 0.00146537f
cc_132 N_NET1_c_188_n N_B_c_252_n 5.75904e-19
cc_133 N_NET1_c_190_n N_B_c_252_n 3.48267e-19
cc_134 N_NET1_c_178_n N_Z_c_256_n 7.69306e-19
*
.ends
*
*
.subckt AND2_HPNW12 A B Y VDD VSS
xgate (VSS VDD A B Y) G3_AND2_N3
.ends
*
* File: G2_AOI21_N3.pex.netlist
* Created: Mon Apr 11 18:50:47 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_AOI21_N3_VSS 2 4 6 8 19 30 35 38 43 48 57 66 67 69 77 78 79 84 86
+ 88 89 Vss
c48 89 Vss 4.28045e-19
c49 86 Vss 0.00576702f
c50 84 Vss 0.00198426f
c51 79 Vss 0.00132518f
c52 78 Vss 4.66086e-19
c53 77 Vss 0.00250771f
c54 69 Vss 0.00104615f
c55 67 Vss 0.0101744f
c56 66 Vss 0.00354326f
c57 65 Vss 0.00133883f
c58 57 Vss 0.00699915f
c59 48 Vss 2.01624e-19
c60 43 Vss 0.00190058f
c61 38 Vss 0.00140655f
c62 35 Vss 0.00813966f
c63 30 Vss 0.0101549f
c64 25 Vss 0.0829032f
c65 19 Vss 0.0350566f
c66 18 Vss 0.0688416f
c67 8 Vss 0.190897f
c68 4 Vss 0.189497f
r69 85 89 0.551426
r70 85 86 18.3386
r71 84 89 0.551426
r72 83 84 5.50157
r73 79 89 0.0828784
r74 77 86 0.652036
r75 77 78 4.33457
r76 73 78 0.652036
r77 68 88 0.326149
r78 67 83 0.652298
r79 67 68 15.1308
r80 66 69 0.655813
r81 65 88 0.326149
r82 65 66 5.50157
r83 48 79 1.82344
r84 43 57 1.16709
r85 43 73 2.16729
r86 38 69 1.82344
r87 35 48 1.16709
r88 30 38 1.16709
r89 25 57 0.0476429
r90 23 25 2.04225
r91 20 23 0.0685365
r92 18 23 0.5835
r93 18 19 2.8008
r94 15 19 0.652036
r95 8 20 5.1348
r96 6 35 0.123773
r97 4 15 5.1348
r98 2 30 0.123773
.ends

.subckt PM_G2_AOI21_N3_VDD 2 4 6 8 10 29 37 42 45 46 48 50 54 56 57 58 63 65 66
+ 68 74 Vss
c56 74 Vss 0.004704f
c57 66 Vss 4.52364e-19
c58 65 Vss 0.00371658f
c59 63 Vss 0.0104139f
c60 58 Vss 0.0017471f
c61 57 Vss 6.04409e-19
c62 56 Vss 0.00309603f
c63 54 Vss 0.00137895f
c64 51 Vss 0.00173381f
c65 50 Vss 0.0117653f
c66 48 Vss 0.00158874f
c67 46 Vss 0.00143356f
c68 45 Vss 0.00419705f
c69 42 Vss 0.0082636f
c70 37 Vss 0.010107f
c71 33 Vss 0.0307825f
c72 29 Vss 8.92604e-20
c73 26 Vss 0.101624f
c74 22 Vss 0.0359157f
c75 21 Vss 0.0712517f
c76 8 Vss 0.189919f
c77 6 Vss 0.190671f
c78 2 Vss 0.189552f
r79 65 68 0.326018
r80 64 66 0.551426
r81 64 65 5.50157
r82 63 66 0.551426
r83 62 63 18.3386
r84 58 66 0.0828784
r85 58 60 1.82344
r86 56 62 0.652036
r87 56 57 4.37625
r88 54 74 1.16709
r89 52 57 0.652036
r90 52 54 2.16729
r91 50 68 0.326018
r92 50 51 15.6711
r93 46 48 1.82344
r94 45 51 0.652036
r95 44 46 0.655813
r96 44 45 5.50157
r97 42 60 1.16709
r98 37 48 1.16709
r99 29 74 0.0476429
r100 27 33 0.494161
r101 27 29 1.45875
r102 26 30 0.652036
r103 26 29 1.45875
r104 23 33 0.128424
r105 21 33 0.494161
r106 21 22 2.8008
r107 18 22 0.652036
r108 10 42 0.123773
r109 8 30 5.1348
r110 6 23 5.1348
r111 4 37 0.123773
r112 2 18 5.1348
.ends

.subckt PM_G2_AOI21_N3_B 2 4 20 23 26 29 Vss
c18 29 Vss 0.00496711f
c19 23 Vss 4.14813e-19
c20 20 Vss 0.0923936f
c21 16 Vss 0.0610957f
c22 4 Vss 0.211686f
c23 2 Vss 0.427124f
r24 23 29 1.16709
r25 23 26 0.125036
r26 18 20 2.04225
r27 16 29 0.197068
r28 13 16 1.2837
r29 10 20 0.0685365
r30 8 18 0.0685365
r31 7 13 0.0685365
r32 4 10 5.6016
r33 2 8 11.2032
r34 2 7 5.1348
.ends

.subckt PM_G2_AOI21_N3_C 2 4 6 17 24 28 31 36 39 43 56 Vss
c47 56 Vss 0.00111429f
c48 43 Vss 0.0052438f
c49 39 Vss 0.00260114f
c50 36 Vss 3.26162e-19
c51 31 Vss 0.00720813f
c52 28 Vss 0.0949366f
c53 24 Vss 0.084323f
c54 17 Vss 4.93054e-19
c55 6 Vss 0.286419f
c56 4 Vss 0.25621f
c57 2 Vss 0.189817f
r58 52 56 0.652036
r59 39 56 5.16814
r60 36 39 0.0833571
r61 31 43 1.16709
r62 31 52 12.2535
r63 26 28 2.04225
r64 24 43 0.0476429
r65 21 24 1.92555
r66 18 28 0.0685365
r67 17 39 1.16709
r68 13 26 0.0685365
r69 13 17 2.8008
r70 10 21 0.0685365
r71 6 18 8.4024
r72 4 17 5.6016
r73 2 10 5.1348
.ends

.subckt PM_G2_AOI21_N3_Z 2 4 6 8 23 27 30 33 Vss
c33 30 Vss 0.00262006f
c34 27 Vss 0.00473513f
c35 23 Vss 0.00644988f
c36 8 Vss 0.00143493f
c37 6 Vss 0.00143493f
r38 33 35 7.5855
r39 30 33 5.2515
r40 27 35 1.16709
r41 23 30 1.16709
r42 8 27 0.123773
r43 6 23 0.123773
r44 4 27 0.123773
r45 2 23 0.123773
.ends

.subckt PM_G2_AOI21_N3_A 2 4 10 11 13 14 15 20 24 29 32 Vss
c32 32 Vss 9.42706e-19
c33 29 Vss 5.87748e-19
c34 24 Vss 1.66175e-19
c35 20 Vss 0.191363f
c36 18 Vss 0.0247918f
c37 15 Vss 0.0322409f
c38 14 Vss 0.0740343f
c39 13 Vss 0.0312529f
c40 11 Vss 0.0324985f
c41 10 Vss 0.122088f
c42 2 Vss 0.292885f
r43 26 32 1.16709
r44 26 29 0.0729375
r45 24 32 0.262036
r46 20 32 0.238214
r47 18 24 0.326018
r48 18 20 0.64185
r49 15 24 2.50905
r50 14 24 0.326018
r51 14 24 0.1167
r52 13 15 0.652036
r53 12 13 1.22535
r54 10 12 0.652036
r55 10 11 3.09255
r56 7 11 0.652036
r57 4 20 5.0181
r58 2 7 8.7525
.ends

.subckt G2_AOI21_N3  VSS VDD B C Z A
*
* A	A
* Z	Z
* C	C
* B	B
* VDD	VDD
* VSS	VSS
XI18.X0 N_Z_XI18.X0_D N_VDD_XI18.X0_PGD N_A_XI18.X0_CG N_B_XI18.X0_PGS
+ N_VSS_XI18.X0_S TIGFET_HPNW12
XI16.X0 N_Z_XI16.X0_D N_VSS_XI16.X0_PGD N_B_XI16.X0_CG N_C_XI16.X0_PGS
+ N_VDD_XI16.X0_S TIGFET_HPNW12
XI19.X0 N_Z_XI19.X0_D N_VDD_XI19.X0_PGD N_C_XI19.X0_CG N_VDD_XI19.X0_PGS
+ N_VSS_XI19.X0_S TIGFET_HPNW12
XI17.X0 N_Z_XI17.X0_D N_VSS_XI17.X0_PGD N_A_XI17.X0_CG N_C_XI17.X0_PGS
+ N_VDD_XI17.X0_S TIGFET_HPNW12
*
x_PM_G2_AOI21_N3_VSS N_VSS_XI18.X0_S N_VSS_XI16.X0_PGD N_VSS_XI19.X0_S
+ N_VSS_XI17.X0_PGD N_VSS_c_3_p N_VSS_c_34_p N_VSS_c_8_p N_VSS_c_2_p N_VSS_c_4_p
+ N_VSS_c_9_p N_VSS_c_5_p N_VSS_c_21_p N_VSS_c_10_p N_VSS_c_1_p N_VSS_c_6_p
+ N_VSS_c_7_p N_VSS_c_12_p N_VSS_c_14_p N_VSS_c_15_p VSS N_VSS_c_16_p Vss
+ PM_G2_AOI21_N3_VSS
x_PM_G2_AOI21_N3_VDD N_VDD_XI18.X0_PGD N_VDD_XI16.X0_S N_VDD_XI19.X0_PGD
+ N_VDD_XI19.X0_PGS N_VDD_XI17.X0_S N_VDD_c_76_p N_VDD_c_90_p N_VDD_c_91_p
+ N_VDD_c_75_p N_VDD_c_49_n N_VDD_c_50_n N_VDD_c_51_n N_VDD_c_70_p N_VDD_c_56_n
+ N_VDD_c_59_n N_VDD_c_60_n N_VDD_c_61_n N_VDD_c_65_n N_VDD_c_68_n VDD
+ N_VDD_c_71_p Vss PM_G2_AOI21_N3_VDD
x_PM_G2_AOI21_N3_B N_B_XI18.X0_PGS N_B_XI16.X0_CG N_B_c_113_p N_B_c_105_n B
+ N_B_c_110_n Vss PM_G2_AOI21_N3_B
x_PM_G2_AOI21_N3_C N_C_XI16.X0_PGS N_C_XI19.X0_CG N_C_XI17.X0_PGS N_C_c_135_n
+ N_C_c_137_n N_C_c_138_n N_C_c_124_n C N_C_c_127_n N_C_c_128_n N_C_c_132_n Vss
+ PM_G2_AOI21_N3_C
x_PM_G2_AOI21_N3_Z N_Z_XI18.X0_D N_Z_XI16.X0_D N_Z_XI19.X0_D N_Z_XI17.X0_D
+ N_Z_c_170_n N_Z_c_180_n N_Z_c_174_n Z Vss PM_G2_AOI21_N3_Z
x_PM_G2_AOI21_N3_A N_A_XI18.X0_CG N_A_XI17.X0_CG N_A_c_203_n N_A_c_213_n
+ N_A_c_214_n N_A_c_204_n N_A_c_215_n N_A_c_221_n N_A_c_205_n A N_A_c_207_n Vss
+ PM_G2_AOI21_N3_A
cc_1 N_VSS_c_1_p N_VDD_c_49_n 3.30468e-19
cc_2 N_VSS_c_2_p N_VDD_c_50_n 4.89405e-19
cc_3 N_VSS_c_3_p N_VDD_c_51_n 0.00126279f
cc_4 N_VSS_c_4_p N_VDD_c_51_n 0.00161703f
cc_5 N_VSS_c_5_p N_VDD_c_51_n 2.26455e-19
cc_6 N_VSS_c_6_p N_VDD_c_51_n 0.00345242f
cc_7 N_VSS_c_7_p N_VDD_c_51_n 0.00169823f
cc_8 N_VSS_c_8_p N_VDD_c_56_n 2.74986e-19
cc_9 N_VSS_c_9_p N_VDD_c_56_n 3.26764e-19
cc_10 N_VSS_c_10_p N_VDD_c_56_n 0.00463433f
cc_11 N_VSS_c_10_p N_VDD_c_59_n 0.00166316f
cc_12 N_VSS_c_12_p N_VDD_c_60_n 4.01154e-19
cc_13 N_VSS_c_9_p N_VDD_c_61_n 0.00187494f
cc_14 N_VSS_c_14_p N_VDD_c_61_n 0.00422386f
cc_15 N_VSS_c_15_p N_VDD_c_61_n 0.00869026f
cc_16 N_VSS_c_16_p N_VDD_c_61_n 9.16632e-19
cc_17 N_VSS_c_4_p N_VDD_c_65_n 4.83895e-19
cc_18 N_VSS_c_6_p N_VDD_c_65_n 0.00105311f
cc_19 N_VSS_c_15_p N_VDD_c_65_n 0.00385589f
cc_20 N_VSS_c_15_p N_VDD_c_68_n 0.00115015f
cc_21 N_VSS_c_21_p N_B_c_105_n 3.69138e-19
cc_22 N_VSS_c_10_p N_B_c_105_n 3.72732e-19
cc_23 N_VSS_XI16.X0_PGD N_C_XI16.X0_PGS 0.00150757f
cc_24 N_VSS_c_4_p N_C_c_124_n 8.90801e-19
cc_25 N_VSS_c_5_p N_C_c_124_n 3.44698e-19
cc_26 N_VSS_c_15_p N_C_c_124_n 0.00209922f
cc_27 N_VSS_c_15_p N_C_c_127_n 5.11302e-19
cc_28 N_VSS_XI16.X0_PGD N_C_c_128_n 3.23173e-19
cc_29 N_VSS_c_3_p N_C_c_128_n 0.00480946f
cc_30 N_VSS_c_4_p N_C_c_128_n 3.44698e-19
cc_31 N_VSS_c_5_p N_C_c_128_n 6.61756e-19
cc_32 N_VSS_c_10_p N_C_c_132_n 0.00205555f
cc_33 N_VSS_c_15_p N_C_c_132_n 3.90377e-19
cc_34 N_VSS_c_34_p N_Z_c_170_n 3.43419e-19
cc_35 N_VSS_c_8_p N_Z_c_170_n 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_c_170_n 3.48267e-19
cc_37 N_VSS_c_9_p N_Z_c_170_n 3.48267e-19
cc_38 N_VSS_c_34_p N_Z_c_174_n 3.48267e-19
cc_39 N_VSS_c_8_p N_Z_c_174_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_174_n 5.71987e-19
cc_41 N_VSS_c_9_p N_Z_c_174_n 5.71987e-19
cc_42 N_VSS_c_10_p N_Z_c_174_n 3.02286e-19
cc_43 N_VSS_c_15_p N_Z_c_174_n 9.87738e-19
cc_44 N_VSS_XI16.X0_PGD N_A_c_203_n 7.5154e-19
cc_45 N_VSS_XI17.X0_PGD N_A_c_204_n 0.00163887f
cc_46 N_VSS_c_5_p N_A_c_205_n 5.05931e-19
cc_47 N_VSS_c_5_p A 2.15082e-19
cc_48 N_VSS_c_4_p N_A_c_207_n 2.15082e-19
cc_49 N_VDD_XI18.X0_PGD N_B_XI18.X0_PGS 0.00174385f
cc_50 N_VDD_c_70_p N_B_c_105_n 6.29947e-19
cc_51 N_VDD_c_71_p N_B_c_105_n 3.48267e-19
cc_52 N_VDD_XI18.X0_PGD N_B_c_110_n 3.23173e-19
cc_53 N_VDD_c_70_p N_B_c_110_n 4.44903e-19
cc_54 N_VDD_c_71_p N_B_c_110_n 6.39485e-19
cc_55 N_VDD_c_75_p N_C_XI16.X0_PGS 3.81609e-19
cc_56 N_VDD_c_76_p N_C_c_135_n 5.33384e-19
cc_57 N_VDD_c_61_n N_C_c_135_n 5.92666e-19
cc_58 N_VDD_c_51_n N_C_c_137_n 3.8746e-19
cc_59 N_VDD_XI19.X0_PGS N_C_c_138_n 8.42974e-19
cc_60 N_VDD_c_61_n N_C_c_138_n 6.25289e-19
cc_61 N_VDD_c_75_p N_C_c_124_n 0.00129723f
cc_62 N_VDD_c_50_n N_C_c_124_n 4.34459e-19
cc_63 N_VDD_c_51_n N_C_c_124_n 0.00204347f
cc_64 N_VDD_c_70_p C 2.77106e-19
cc_65 N_VDD_c_61_n C 4.49702e-19
cc_66 N_VDD_c_71_p C 2.15082e-19
cc_67 N_VDD_c_51_n N_C_c_127_n 5.0979e-19
cc_68 N_VDD_c_75_p N_C_c_128_n 3.66936e-19
cc_69 N_VDD_c_51_n N_C_c_128_n 2.64932e-19
cc_70 N_VDD_c_90_p N_Z_c_180_n 3.43419e-19
cc_71 N_VDD_c_91_p N_Z_c_180_n 3.43419e-19
cc_72 N_VDD_c_50_n N_Z_c_180_n 3.72199e-19
cc_73 N_VDD_c_51_n N_Z_c_180_n 2.74986e-19
cc_74 N_VDD_c_60_n N_Z_c_180_n 3.72199e-19
cc_75 N_VDD_c_90_p N_Z_c_174_n 3.48267e-19
cc_76 N_VDD_c_91_p N_Z_c_174_n 3.48267e-19
cc_77 N_VDD_c_50_n N_Z_c_174_n 5.09542e-19
cc_78 N_VDD_c_51_n N_Z_c_174_n 5.72568e-19
cc_79 N_VDD_c_60_n N_Z_c_174_n 7.72285e-19
cc_80 N_VDD_c_61_n N_Z_c_174_n 0.00179861f
cc_81 N_VDD_XI18.X0_PGD N_A_c_203_n 6.25166e-19
cc_82 N_VDD_XI19.X0_PGD N_A_c_204_n 3.70201e-19
cc_83 N_VDD_c_61_n A 4.8807e-19
cc_84 N_VDD_c_61_n N_A_c_207_n 3.66936e-19
cc_85 N_B_c_113_p N_C_XI16.X0_PGS 0.0020206f
cc_86 N_B_XI18.X0_PGS N_C_XI19.X0_CG 2.46172e-19
cc_87 N_B_c_113_p N_C_XI17.X0_PGS 4.66827e-19
cc_88 N_B_c_105_n N_C_c_132_n 2.19701e-19
cc_89 N_B_XI18.X0_PGS N_Z_c_174_n 2.61881e-19
cc_90 N_B_XI18.X0_PGS N_A_XI18.X0_CG 0.00881601f
cc_91 N_B_c_113_p N_A_c_213_n 0.00191565f
cc_92 N_B_XI18.X0_PGS N_A_c_214_n 6.07734e-19
cc_93 N_B_c_113_p N_A_c_215_n 0.00136534f
cc_94 N_B_c_113_p N_A_c_207_n 2.87722e-19
cc_95 N_C_c_135_n N_Z_c_174_n 9.83688e-19
cc_96 N_C_c_124_n N_Z_c_174_n 0.00308891f
cc_97 C N_Z_c_174_n 0.00140888f
cc_98 N_C_c_127_n N_Z_c_174_n 0.00195497f
cc_99 N_C_c_132_n N_Z_c_174_n 2.70867e-19
cc_100 N_C_XI19.X0_CG N_A_XI18.X0_CG 5.48933e-19
cc_101 N_C_c_135_n N_A_XI18.X0_CG 5.60239e-19
cc_102 N_C_XI17.X0_PGS N_A_c_203_n 8.10159e-19
cc_103 N_C_c_138_n N_A_c_203_n 0.00121323f
cc_104 N_C_XI17.X0_PGS N_A_c_221_n 4.42555e-19
cc_105 N_C_c_135_n N_A_c_205_n 9.47282e-19
cc_106 N_C_c_135_n A 4.56568e-19
cc_107 C A 6.3743e-19
cc_108 N_C_XI17.X0_PGS N_A_c_207_n 0.00570455f
cc_109 N_C_c_135_n N_A_c_207_n 6.1245e-19
cc_110 N_C_c_138_n N_A_c_207_n 0.00239404f
cc_111 C N_A_c_207_n 4.56568e-19
cc_112 N_Z_c_174_n N_A_XI18.X0_CG 5.52516e-19
cc_113 N_Z_c_170_n N_A_c_203_n 3.56294e-19
cc_114 N_Z_c_174_n N_A_c_203_n 3.092e-19
cc_115 N_Z_c_180_n N_A_c_215_n 5.66216e-19
cc_116 N_Z_c_174_n A 0.00149422f
cc_117 N_Z_c_174_n N_A_c_207_n 9.53426e-19
*
.ends
*
*
.subckt AOI21_HPNW12 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 B0 Y A0) G2_AOI21_N3
.ends
*
* File: G2_BUF1_N3.pex.netlist
* Created: Wed Mar  2 15:50:41 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_BUF1_N3_VDD 2 4 7 11 28 30 32 44 48 52 54 56 57 61 65 67 71 75 78
+ 90 95 Vss
c55 95 Vss 0.00494983f
c56 90 Vss 0.00475556f
c57 80 Vss 9.22237e-19
c58 79 Vss 9.22237e-19
c59 75 Vss 0.00138508f
c60 71 Vss 9.81533e-19
c61 68 Vss 0.00177515f
c62 67 Vss 0.00751016f
c63 65 Vss 0.0012592f
c64 61 Vss 0.0012592f
c65 57 Vss 0.00744668f
c66 56 Vss 0.00466777f
c67 54 Vss 0.00779694f
c68 52 Vss 0.00466777f
c69 51 Vss 0.00177515f
c70 48 Vss 0.00810125f
c71 44 Vss 0.0100206f
c72 32 Vss 0.0356247f
c73 31 Vss 0.102427f
c74 28 Vss 0.0356247f
c75 27 Vss 0.102427f
c76 11 Vss 0.378484f
c77 7 Vss 0.378484f
r78 75 95 1.16709
r79 73 75 2.16729
r80 71 90 1.16709
r81 69 71 2.16729
r82 67 73 0.652036
r83 67 68 10.1279
r84 63 80 0.0828784
r85 63 65 1.82344
r86 59 79 0.0828784
r87 59 61 1.82344
r88 58 78 0.326018
r89 57 69 0.652036
r90 57 58 10.1279
r91 56 68 0.652036
r92 55 80 0.551426
r93 55 56 5.50157
r94 54 80 0.551426
r95 53 79 0.551426
r96 53 54 8.58579
r97 52 79 0.551426
r98 51 78 0.326018
r99 51 52 5.50157
r100 48 65 1.16709
r101 44 61 1.16709
r102 34 95 0.0476429
r103 32 34 1.45875
r104 31 38 0.652036
r105 31 34 1.45875
r106 30 90 0.0476429
r107 28 30 1.45875
r108 27 35 0.652036
r109 27 30 1.45875
r110 24 32 0.652036
r111 21 28 0.652036
r112 11 38 5.1348
r113 11 24 5.1348
r114 7 35 5.1348
r115 7 21 5.1348
r116 4 48 0.123773
r117 2 44 0.123773
.ends

.subckt PM_G2_BUF1_N3_VSS 3 7 10 12 27 28 31 32 45 49 52 57 62 67 72 77 97 98 99
+ 100 101 105 110 112 114 116 Vss
c52 118 Vss 6.78504e-19
c53 117 Vss 6.78504e-19
c54 114 Vss 0.00360796f
c55 112 Vss 0.00582053f
c56 110 Vss 0.00360796f
c57 109 Vss 0.0013648f
c58 105 Vss 0.0010737f
c59 101 Vss 9.14356e-19
c60 100 Vss 5.83649e-19
c61 99 Vss 0.00682958f
c62 98 Vss 5.83649e-19
c63 97 Vss 0.00550031f
c64 77 Vss 0.00392669f
c65 72 Vss 0.00392498f
c66 67 Vss 1.62518e-19
c67 62 Vss 7.10513e-22
c68 57 Vss 8.49747e-19
c69 52 Vss 0.00100529f
c70 49 Vss 0.0100686f
c71 45 Vss 0.00814922f
c72 32 Vss 0.0350852f
c73 31 Vss 0.0994129f
c74 28 Vss 0.0350852f
c75 27 Vss 0.0994129f
c76 7 Vss 0.377694f
c77 3 Vss 0.377694f
r78 113 118 0.551426
r79 113 114 5.50157
r80 112 118 0.551426
r81 111 117 0.551426
r82 111 112 8.58579
r83 110 117 0.551426
r84 109 116 0.326018
r85 109 110 5.50157
r86 105 118 0.0828784
r87 101 117 0.0828784
r88 99 114 0.652036
r89 99 100 10.1279
r90 97 116 0.326018
r91 97 98 10.1279
r92 93 100 0.652036
r93 89 98 0.652036
r94 67 105 1.82344
r95 62 101 1.82344
r96 57 77 1.16709
r97 57 93 2.16729
r98 52 72 1.16709
r99 52 89 2.16729
r100 49 67 1.16709
r101 45 62 1.16709
r102 34 77 0.0476429
r103 32 34 1.45875
r104 31 38 0.652036
r105 31 34 1.45875
r106 30 72 0.0476429
r107 28 30 1.45875
r108 27 35 0.652036
r109 27 30 1.45875
r110 24 32 0.652036
r111 21 28 0.652036
r112 12 49 0.123773
r113 10 45 0.123773
r114 7 38 5.1348
r115 7 24 5.1348
r116 3 35 5.1348
r117 3 21 5.1348
.ends

.subckt PM_G2_BUF1_N3_A 2 4 12 24 27 Vss
c13 27 Vss 0.00315166f
c14 24 Vss 1.56823e-19
c15 12 Vss 0.20431f
c16 9 Vss 0.180512f
c17 7 Vss 0.0247918f
c18 4 Vss 0.193588f
r19 24 27 1.16709
r20 15 27 0.0476429
r21 13 15 0.326018
r22 13 15 0.1167
r23 12 16 0.652036
r24 12 15 6.7686
r25 9 27 0.357321
r26 7 15 0.326018
r27 7 9 0.40845
r28 4 16 5.1348
r29 2 9 4.72635
.ends

.subckt PM_G2_BUF1_N3_Z 2 4 13 16 19 Vss
c13 16 Vss 3.73795e-19
c14 13 Vss 0.00513911f
c15 4 Vss 0.00176592f
r16 16 19 0.0416786
r17 13 16 1.16709
r18 4 13 0.123773
r19 2 13 0.123773
.ends

.subckt PM_G2_BUF1_N3_NET17 2 4 6 8 18 33 36 41 50 58 Vss
c31 58 Vss 5.10694e-19
c32 50 Vss 0.0034988f
c33 41 Vss 0.0021514f
c34 36 Vss 0.0018043f
c35 33 Vss 0.00513911f
c36 22 Vss 0.0247918f
c37 19 Vss 0.0299669f
c38 18 Vss 0.173331f
c39 8 Vss 0.00176592f
c40 6 Vss 0.180667f
c41 2 Vss 0.192541f
r42 54 58 0.653045
r43 41 50 1.16709
r44 41 58 2.1395
r45 36 54 5.29318
r46 33 36 1.16709
r47 28 50 0.0476429
r48 26 50 0.357321
r49 22 28 0.326018
r50 22 26 0.40845
r51 19 28 6.7686
r52 18 28 0.326018
r53 18 28 0.1167
r54 15 19 0.652036
r55 8 33 0.123773
r56 6 26 4.72635
r57 4 33 0.123773
r58 2 15 5.1348
.ends

.subckt G2_BUF1_N3  VDD VSS A Z
*
* Z	Z
* A	A
* VSS	VSS
* VDD	VDD
XI14.X0 N_Z_XI14.X0_D N_VSS_XI14.X0_PGD N_NET17_XI14.X0_CG N_VSS_XI14.X0_PGD
+ N_VDD_XI14.X0_S TIGFET_HPNW12
XI11.X0 N_NET17_XI11.X0_D N_VSS_XI11.X0_PGD N_A_XI11.X0_CG N_VSS_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW12
XI13.X0 N_Z_XI13.X0_D N_VDD_XI13.X0_PGD N_NET17_XI13.X0_CG N_VDD_XI13.X0_PGD
+ N_VSS_XI13.X0_S TIGFET_HPNW12
XI12.X0 N_NET17_XI12.X0_D N_VDD_XI12.X0_PGD N_A_XI12.X0_CG N_VDD_XI12.X0_PGD
+ N_VSS_XI12.X0_S TIGFET_HPNW12
*
x_PM_G2_BUF1_N3_VDD N_VDD_XI14.X0_S N_VDD_XI11.X0_S N_VDD_XI13.X0_PGD
+ N_VDD_XI12.X0_PGD N_VDD_c_4_p N_VDD_c_50_p N_VDD_c_8_p N_VDD_c_36_p
+ N_VDD_c_45_p N_VDD_c_6_p N_VDD_c_34_p N_VDD_c_3_p N_VDD_c_5_p N_VDD_c_38_p
+ N_VDD_c_46_p N_VDD_c_9_p N_VDD_c_13_p N_VDD_c_17_p VDD N_VDD_c_14_p
+ N_VDD_c_18_p Vss PM_G2_BUF1_N3_VDD
x_PM_G2_BUF1_N3_VSS N_VSS_XI14.X0_PGD N_VSS_XI11.X0_PGD N_VSS_XI13.X0_S
+ N_VSS_XI12.X0_S N_VSS_c_59_n N_VSS_c_61_n N_VSS_c_63_n N_VSS_c_65_n
+ N_VSS_c_93_p N_VSS_c_99_p N_VSS_c_66_n N_VSS_c_70_n N_VSS_c_94_p N_VSS_c_100_p
+ N_VSS_c_74_n N_VSS_c_78_n N_VSS_c_81_n N_VSS_c_82_n N_VSS_c_83_n N_VSS_c_84_n
+ N_VSS_c_96_p N_VSS_c_103_p N_VSS_c_85_n N_VSS_c_104_p N_VSS_c_86_n VSS Vss
+ PM_G2_BUF1_N3_VSS
x_PM_G2_BUF1_N3_A N_A_XI11.X0_CG N_A_XI12.X0_CG N_A_c_108_n A N_A_c_111_n Vss
+ PM_G2_BUF1_N3_A
x_PM_G2_BUF1_N3_Z N_Z_XI14.X0_D N_Z_XI13.X0_D N_Z_c_121_n N_Z_c_124_n Z Vss
+ PM_G2_BUF1_N3_Z
x_PM_G2_BUF1_N3_NET17 N_NET17_XI14.X0_CG N_NET17_XI11.X0_D N_NET17_XI13.X0_CG
+ N_NET17_XI12.X0_D N_NET17_c_135_n N_NET17_c_137_n N_NET17_c_139_n
+ N_NET17_c_142_n N_NET17_c_146_n N_NET17_c_147_n Vss PM_G2_BUF1_N3_NET17
cc_1 N_VDD_XI13.X0_PGD N_VSS_XI14.X0_PGD 0.00200662f
cc_2 N_VDD_XI12.X0_PGD N_VSS_XI11.X0_PGD 0.00200662f
cc_3 N_VDD_c_3_p N_VSS_XI11.X0_PGD 4.00543e-19
cc_4 N_VDD_c_4_p N_VSS_c_59_n 0.00200662f
cc_5 N_VDD_c_5_p N_VSS_c_59_n 3.89167e-19
cc_6 N_VDD_c_6_p N_VSS_c_61_n 4.00543e-19
cc_7 N_VDD_c_5_p N_VSS_c_61_n 4.0633e-19
cc_8 N_VDD_c_8_p N_VSS_c_63_n 0.00200662f
cc_9 N_VDD_c_9_p N_VSS_c_63_n 3.89167e-19
cc_10 N_VDD_c_9_p N_VSS_c_65_n 4.0633e-19
cc_11 N_VDD_c_6_p N_VSS_c_66_n 9.94764e-19
cc_12 N_VDD_c_5_p N_VSS_c_66_n 0.00162079f
cc_13 N_VDD_c_13_p N_VSS_c_66_n 0.00106273f
cc_14 N_VDD_c_14_p N_VSS_c_66_n 3.48267e-19
cc_15 N_VDD_c_3_p N_VSS_c_70_n 9.94764e-19
cc_16 N_VDD_c_9_p N_VSS_c_70_n 0.00141604f
cc_17 N_VDD_c_17_p N_VSS_c_70_n 0.00110056f
cc_18 N_VDD_c_18_p N_VSS_c_70_n 3.48267e-19
cc_19 N_VDD_c_6_p N_VSS_c_74_n 3.66936e-19
cc_20 N_VDD_c_5_p N_VSS_c_74_n 2.2543e-19
cc_21 N_VDD_c_13_p N_VSS_c_74_n 3.99794e-19
cc_22 N_VDD_c_14_p N_VSS_c_74_n 6.489e-19
cc_23 N_VDD_c_3_p N_VSS_c_78_n 3.66936e-19
cc_24 N_VDD_c_9_p N_VSS_c_78_n 0.00114409f
cc_25 N_VDD_c_18_p N_VSS_c_78_n 6.489e-19
cc_26 N_VDD_c_5_p N_VSS_c_81_n 0.00589548f
cc_27 N_VDD_c_5_p N_VSS_c_82_n 0.0017359f
cc_28 N_VDD_c_9_p N_VSS_c_83_n 0.00593021f
cc_29 N_VDD_c_9_p N_VSS_c_84_n 0.0017359f
cc_30 N_VDD_c_13_p N_VSS_c_85_n 3.85245e-19
cc_31 N_VDD_c_17_p N_VSS_c_86_n 3.85245e-19
cc_32 N_VDD_XI13.X0_PGD N_A_c_108_n 4.14544e-19
cc_33 N_VDD_XI12.X0_PGD N_A_c_108_n 4.09718e-19
cc_34 N_VDD_c_34_p A 9.3432e-19
cc_35 N_VDD_c_34_p N_A_c_111_n 5.79991e-19
cc_36 N_VDD_c_36_p N_Z_c_121_n 3.43419e-19
cc_37 N_VDD_c_5_p N_Z_c_121_n 2.74986e-19
cc_38 N_VDD_c_38_p N_Z_c_121_n 3.72199e-19
cc_39 N_VDD_c_36_p N_Z_c_124_n 3.48267e-19
cc_40 N_VDD_c_5_p N_Z_c_124_n 3.66281e-19
cc_41 N_VDD_c_38_p N_Z_c_124_n 7.4527e-19
cc_42 N_VDD_c_34_p N_NET17_XI14.X0_CG 3.93898e-19
cc_43 N_VDD_XI13.X0_PGD N_NET17_c_135_n 4.09718e-19
cc_44 N_VDD_XI12.X0_PGD N_NET17_c_135_n 4.14544e-19
cc_45 N_VDD_c_45_p N_NET17_c_137_n 3.43419e-19
cc_46 N_VDD_c_46_p N_NET17_c_137_n 3.72199e-19
cc_47 N_VDD_c_45_p N_NET17_c_139_n 3.48267e-19
cc_48 N_VDD_c_46_p N_NET17_c_139_n 8.0086e-19
cc_49 N_VDD_c_9_p N_NET17_c_139_n 3.21336e-19
cc_50 N_VDD_c_50_p N_NET17_c_142_n 2.21762e-19
cc_51 N_VDD_c_34_p N_NET17_c_142_n 2.74452e-19
cc_52 N_VDD_c_13_p N_NET17_c_142_n 2.88301e-19
cc_53 N_VDD_c_14_p N_NET17_c_142_n 2.30774e-19
cc_54 N_VDD_c_13_p N_NET17_c_146_n 2.28697e-19
cc_55 N_VDD_c_34_p N_NET17_c_147_n 7.45369e-19
cc_56 N_VSS_XI14.X0_PGD N_A_c_108_n 4.14544e-19
cc_57 N_VSS_XI11.X0_PGD N_A_c_108_n 4.09718e-19
cc_58 N_VSS_c_66_n A 2.26871e-19
cc_59 N_VSS_c_70_n A 3.35067e-19
cc_60 N_VSS_c_78_n A 2.30774e-19
cc_61 N_VSS_c_70_n N_A_c_111_n 2.28892e-19
cc_62 N_VSS_c_93_p N_Z_c_121_n 3.43419e-19
cc_63 N_VSS_c_94_p N_Z_c_121_n 3.48267e-19
cc_64 N_VSS_c_94_p N_Z_c_124_n 5.37696e-19
cc_65 N_VSS_c_96_p N_Z_c_124_n 2.7826e-19
cc_66 N_VSS_XI14.X0_PGD N_NET17_c_135_n 4.09718e-19
cc_67 N_VSS_XI11.X0_PGD N_NET17_c_135_n 4.14544e-19
cc_68 N_VSS_c_99_p N_NET17_c_137_n 3.43419e-19
cc_69 N_VSS_c_100_p N_NET17_c_137_n 3.48267e-19
cc_70 N_VSS_c_100_p N_NET17_c_139_n 4.8288e-19
cc_71 N_VSS_c_83_n N_NET17_c_139_n 3.94979e-19
cc_72 N_VSS_c_103_p N_NET17_c_139_n 5.49885e-19
cc_73 N_VSS_c_104_p N_NET17_c_139_n 0.00142716f
cc_74 N_VSS_c_104_p N_NET17_c_142_n 0.00119345f
cc_75 N_VSS_c_81_n N_NET17_c_147_n 6.75516e-19
cc_76 N_VSS_c_83_n N_NET17_c_147_n 4.01006e-19
cc_77 N_A_c_108_n N_NET17_c_135_n 0.00945061f
cc_78 N_A_c_108_n N_NET17_c_137_n 4.98287e-19
cc_79 A N_NET17_c_139_n 8.54729e-19
cc_80 N_Z_c_121_n N_NET17_c_135_n 4.98287e-19
cc_81 N_Z_c_121_n N_NET17_c_137_n 3.80999e-19
cc_82 N_Z_c_124_n N_NET17_c_147_n 2.07279e-19
*
.ends
*
*
.subckt BUF1_HPNW12 A Y VDD VSS
xgate (VDD VSS A Y) G2_BUF1_N3
.ends
*
* File: G3_DFFQ1_N3.pex.netlist
* Created: Wed Apr  6 11:25:19 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_DFFQ1_N3_VSS 2 4 6 8 10 12 14 29 42 44 49 55 59 64 67 72 78 83 88
+ 93 102 111 117 126 127 128 129 133 138 143 149 155 157 162 164 166 167 168 Vss
c101 168 Vss 4.28045e-19
c102 167 Vss 3.75522e-19
c103 166 Vss 3.75522e-19
c104 165 Vss 6.20041e-19
c105 164 Vss 0.00614697f
c106 162 Vss 0.00220014f
c107 157 Vss 0.0014078f
c108 155 Vss 0.00256807f
c109 149 Vss 0.00450029f
c110 143 Vss 0.00309494f
c111 133 Vss 0.00200475f
c112 129 Vss 6.50617e-19
c113 128 Vss 8.16747e-19
c114 127 Vss 0.00572724f
c115 126 Vss 0.0020774f
c116 117 Vss 0.00492488f
c117 111 Vss 0.00403629f
c118 102 Vss 0.00419844f
c119 93 Vss 2.01624e-19
c120 88 Vss 9.8978e-19
c121 83 Vss 8.45647e-19
c122 78 Vss 0.00151704f
c123 72 Vss 0.0130885f
c124 67 Vss 0.00136241f
c125 64 Vss 0.0111802f
c126 59 Vss 0.00964026f
c127 55 Vss 0.00801889f
c128 49 Vss 0.0568987f
c129 44 Vss 0.0568992f
c130 42 Vss 8.92801e-20
c131 29 Vss 0.0356247f
c132 28 Vss 0.101312f
c133 14 Vss 0.189842f
c134 8 Vss 0.191315f
c135 6 Vss 0.188337f
c136 4 Vss 0.188444f
r137 163 168 0.551426
r138 163 164 18.3386
r139 162 168 0.551426
r140 161 162 5.54325
r141 157 168 0.0828784
r142 156 167 0.494161
r143 155 164 0.652036
r144 155 156 4.37625
r145 151 167 0.128424
r146 150 166 0.494161
r147 149 161 0.652036
r148 149 150 10.1279
r149 145 166 0.128424
r150 144 165 0.494161
r151 143 167 0.494161
r152 143 144 7.46046
r153 139 165 0.128424
r154 133 165 0.494161
r155 133 138 1.00029
r156 127 166 0.494161
r157 127 128 15.8795
r158 126 129 0.655813
r159 125 128 0.652036
r160 125 126 5.54325
r161 111 114 0.05
r162 93 157 1.82344
r163 88 117 1.16709
r164 88 151 2.16729
r165 83 114 1.16709
r166 83 145 2.20896
r167 78 139 6.16843
r168 75 138 1.29204
r169 72 102 1.16709
r170 72 75 15.5878
r171 67 129 1.82344
r172 64 93 1.16709
r173 59 78 1.16709
r174 55 67 1.16709
r175 49 117 0.197068
r176 46 49 1.2837
r177 42 111 0.197068
r178 42 44 1.2837
r179 38 46 0.0685365
r180 35 44 0.0685365
r181 31 102 0.0476429
r182 29 31 1.45875
r183 28 32 0.652036
r184 28 31 1.45875
r185 25 29 0.652036
r186 14 38 5.1348
r187 12 64 0.123773
r188 10 59 0.123773
r189 8 35 5.1348
r190 6 32 5.1348
r191 4 25 5.1348
r192 2 55 0.123773
.ends

.subckt PM_G3_DFFQ1_N3_CK 2 4 6 8 18 21 25 35 41 Vss
c33 41 Vss 0.00492267f
c34 35 Vss 3.25681e-19
c35 33 Vss 0.0299314f
c36 25 Vss 0.166167f
c37 21 Vss 8.92801e-20
c38 18 Vss 0.18663f
c39 15 Vss 0.180502f
c40 13 Vss 0.0247918f
c41 6 Vss 0.659388f
c42 4 Vss 0.191169f
r43 41 44 0.05
r44 38 44 1.16709
r45 35 38 0.0416786
r46 26 33 0.494161
r47 25 27 0.652036
r48 25 26 4.84305
r49 22 33 0.128424
r50 21 41 0.0238214
r51 19 21 0.326018
r52 19 21 0.1167
r53 18 33 0.494161
r54 18 21 6.7686
r55 15 41 0.357321
r56 13 21 0.326018
r57 13 15 0.3501
r58 6 8 17.9718
r59 6 27 5.1348
r60 4 22 5.1348
r61 2 15 4.7847
.ends

.subckt PM_G3_DFFQ1_N3_VDD 2 4 6 8 10 12 14 28 42 44 49 56 60 63 64 65 70 72 76
+ 78 79 82 84 86 91 93 95 96 98 99 100 102 104 113 118 Vss
c107 118 Vss 0.00533757f
c108 113 Vss 0.00573314f
c109 104 Vss 0.00489453f
c110 100 Vss 4.52364e-19
c111 99 Vss 2.39889e-19
c112 98 Vss 4.43992e-19
c113 96 Vss 0.00375805f
c114 95 Vss 4.90076e-19
c115 93 Vss 0.00385631f
c116 91 Vss 0.0108071f
c117 86 Vss 0.00177107f
c118 84 Vss 0.0031515f
c119 82 Vss 0.00100814f
c120 79 Vss 4.90412e-19
c121 78 Vss 0.00546064f
c122 76 Vss 6.46297e-19
c123 72 Vss 0.00354521f
c124 70 Vss 0.00226527f
c125 67 Vss 0.00183337f
c126 65 Vss 8.65196e-19
c127 64 Vss 0.00754197f
c128 63 Vss 0.00697044f
c129 60 Vss 0.0112146f
c130 56 Vss 0.0070753f
c131 49 Vss 0.0589116f
c132 44 Vss 0.0581535f
c133 42 Vss 7.85965e-20
c134 29 Vss 0.0372509f
c135 28 Vss 0.101007f
c136 12 Vss 0.191734f
c137 10 Vss 0.189852f
c138 8 Vss 0.00143493f
c139 4 Vss 0.190684f
c140 2 Vss 0.189513f
r141 118 121 0.05
r142 95 104 1.16709
r143 95 96 0.470345
r144 93 102 0.326018
r145 92 100 0.551426
r146 92 93 5.50157
r147 91 100 0.551426
r148 90 91 18.3803
r149 86 100 0.0828784
r150 86 88 1.82344
r151 85 99 0.494161
r152 84 90 0.652036
r153 84 85 4.37625
r154 82 121 1.16709
r155 80 99 0.128424
r156 80 82 2.20896
r157 78 102 0.326018
r158 78 79 10.1279
r159 76 113 1.16709
r160 74 79 0.652036
r161 74 76 2.16729
r162 73 98 0.494161
r163 72 99 0.494161
r164 72 73 7.46046
r165 68 98 0.128424
r166 68 70 6.21011
r167 67 96 3.82922
r168 64 98 0.494161
r169 64 65 13.0037
r170 63 67 0.655813
r171 62 65 0.652036
r172 62 63 10.2113
r173 60 88 1.16709
r174 56 70 1.16709
r175 49 118 0.197068
r176 46 49 1.2837
r177 42 113 0.197068
r178 42 44 1.2837
r179 38 46 0.0685365
r180 35 44 0.0685365
r181 31 104 0.0476429
r182 29 31 1.45875
r183 28 32 0.652036
r184 28 31 1.45875
r185 25 29 0.652036
r186 14 60 0.123773
r187 12 38 5.1348
r188 10 35 5.1348
r189 8 56 0.123773
r190 6 56 0.123773
r191 4 25 5.1348
r192 2 32 5.1348
.ends

.subckt PM_G3_DFFQ1_N3_CKN 2 4 6 8 18 25 28 33 50 Vss
c37 51 Vss 0.00128789f
c38 50 Vss 0.00701318f
c39 33 Vss 3.33899e-19
c40 28 Vss 0.00179767f
c41 25 Vss 0.00520172f
c42 18 Vss 7.22113e-19
c43 6 Vss 0.584002f
c44 4 Vss 0.00143493f
r45 50 51 14.6709
r46 46 51 0.652036
r47 33 50 0.531835
r48 28 46 5.835
r49 25 28 1.16709
r50 18 33 1.16709
r51 8 18 8.9859
r52 6 18 8.9859
r53 4 25 0.123773
r54 2 25 0.123773
.ends

.subckt PM_G3_DFFQ1_N3_D 2 4 11 12 22 25 28 Vss
c24 28 Vss 0.00196994f
c25 25 Vss 4.67436e-19
c26 12 Vss 0.214507f
c27 11 Vss 8.44702e-20
c28 7 Vss 0.0247918f
c29 4 Vss 0.191884f
c30 2 Vss 0.180391f
r31 25 28 1.16709
r32 22 25 0.0364688
r33 15 28 0.0476429
r34 13 15 0.326018
r35 13 15 0.1167
r36 12 16 0.652036
r37 12 15 6.7686
r38 11 28 0.357321
r39 7 15 0.326018
r40 7 11 0.40845
r41 4 16 5.1348
r42 2 11 4.72635
.ends

.subckt PM_G3_DFFQ1_N3_X 2 4 6 8 17 20 23 33 35 39 41 47 Vss
c46 47 Vss 0.00165819f
c47 41 Vss 5.1586e-19
c48 39 Vss 0.00126373f
c49 35 Vss 0.00198822f
c50 33 Vss 0.00525025f
c51 23 Vss 7.81442e-20
c52 20 Vss 0.214848f
c53 17 Vss 0.180344f
c54 15 Vss 0.0247918f
c55 8 Vss 0.191809f
c56 6 Vss 0.00143493f
r57 44 47 1.16709
r58 41 44 2.08393
r59 37 39 6.16843
r60 36 41 0.0685365
r61 35 37 0.652036
r62 35 36 1.70882
r63 33 39 1.16709
r64 23 47 0.0476429
r65 21 23 0.326018
r66 21 23 0.1167
r67 20 24 0.652036
r68 20 23 6.7686
r69 17 47 0.357321
r70 15 23 0.326018
r71 15 17 0.40845
r72 8 24 5.1348
r73 6 33 0.123773
r74 4 17 4.72635
r75 2 33 0.123773
.ends

.subckt PM_G3_DFFQ1_N3_Q 2 4 13 16 Vss
c12 16 Vss 3.46649e-19
c13 13 Vss 0.0045421f
c14 4 Vss 0.00143493f
r15 16 19 0.0416786
r16 13 19 1.16709
r17 4 13 0.123773
r18 2 13 0.123773
.ends

.subckt G3_DFFQ1_N3  VSS CK VDD D Q
*
* Q	Q
* D	D
* VDD	VDD
* CK	CK
* VSS	VSS
XI0.X0 N_CKN_XI0.X0_D N_VDD_XI0.X0_PGD N_CK_XI0.X0_CG N_VDD_XI0.X0_PGS
+ N_VSS_XI0.X0_S TIGFET_HPNW12
XI1.X0 N_CKN_XI1.X0_D N_VSS_XI1.X0_PGD N_CK_XI1.X0_CG N_VSS_XI1.X0_PGS
+ N_VDD_XI1.X0_S TIGFET_HPNW12
XI13.X0 N_X_XI13.X0_D N_VSS_XI13.X0_PGD N_D_XI13.X0_CG N_CK_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW12
XI4.X0 N_Q_XI4.X0_D N_VDD_XI4.X0_PGD N_X_XI4.X0_CG N_CK_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW12
XI12.X0 N_X_XI12.X0_D N_VDD_XI12.X0_PGD N_D_XI12.X0_CG N_CKN_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW12
XI5.X0 N_Q_XI5.X0_D N_VSS_XI5.X0_PGD N_X_XI5.X0_CG N_CKN_XI5.X0_PGS
+ N_VDD_XI5.X0_S TIGFET_HPNW12
*
x_PM_G3_DFFQ1_N3_VSS N_VSS_XI0.X0_S N_VSS_XI1.X0_PGD N_VSS_XI1.X0_PGS
+ N_VSS_XI13.X0_PGD N_VSS_XI4.X0_S N_VSS_XI12.X0_S N_VSS_XI5.X0_PGD N_VSS_c_11_p
+ N_VSS_c_81_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_14_p N_VSS_c_99_p N_VSS_c_41_p
+ N_VSS_c_15_p N_VSS_c_3_p N_VSS_c_30_p N_VSS_c_21_p N_VSS_c_31_p N_VSS_c_42_p
+ N_VSS_c_54_p N_VSS_c_4_p N_VSS_c_34_p N_VSS_c_16_p N_VSS_c_7_p N_VSS_c_20_p
+ N_VSS_c_17_p N_VSS_c_78_p VSS N_VSS_c_35_p N_VSS_c_27_p N_VSS_c_36_p
+ N_VSS_c_44_p N_VSS_c_46_p N_VSS_c_47_p N_VSS_c_28_p N_VSS_c_37_p N_VSS_c_48_p
+ Vss PM_G3_DFFQ1_N3_VSS
x_PM_G3_DFFQ1_N3_CK N_CK_XI0.X0_CG N_CK_XI1.X0_CG N_CK_XI13.X0_PGS
+ N_CK_XI4.X0_PGS N_CK_c_106_n N_CK_c_124_p N_CK_c_107_n CK N_CK_c_114_p Vss
+ PM_G3_DFFQ1_N3_CK
x_PM_G3_DFFQ1_N3_VDD N_VDD_XI0.X0_PGD N_VDD_XI0.X0_PGS N_VDD_XI1.X0_S
+ N_VDD_XI13.X0_S N_VDD_XI4.X0_PGD N_VDD_XI12.X0_PGD N_VDD_XI5.X0_S
+ N_VDD_c_138_n N_VDD_c_224_p N_VDD_c_139_n N_VDD_c_140_n N_VDD_c_197_n
+ N_VDD_c_236_p N_VDD_c_141_n N_VDD_c_145_n N_VDD_c_147_n N_VDD_c_148_n
+ N_VDD_c_150_n N_VDD_c_156_n N_VDD_c_159_n N_VDD_c_165_n N_VDD_c_166_n
+ N_VDD_c_168_n N_VDD_c_171_n N_VDD_c_172_n N_VDD_c_176_n N_VDD_c_180_n
+ N_VDD_c_182_n N_VDD_c_184_n N_VDD_c_185_n N_VDD_c_186_n VDD N_VDD_c_187_n
+ N_VDD_c_189_n N_VDD_c_192_n Vss PM_G3_DFFQ1_N3_VDD
x_PM_G3_DFFQ1_N3_CKN N_CKN_XI0.X0_D N_CKN_XI1.X0_D N_CKN_XI12.X0_PGS
+ N_CKN_XI5.X0_PGS N_CKN_c_257_n N_CKN_c_242_n N_CKN_c_244_n N_CKN_c_248_n
+ N_CKN_c_249_n Vss PM_G3_DFFQ1_N3_CKN
x_PM_G3_DFFQ1_N3_D N_D_XI13.X0_CG N_D_XI12.X0_CG N_D_c_279_n N_D_c_280_n D
+ N_D_c_281_n N_D_c_284_n Vss PM_G3_DFFQ1_N3_D
x_PM_G3_DFFQ1_N3_X N_X_XI13.X0_D N_X_XI4.X0_CG N_X_XI12.X0_D N_X_XI5.X0_CG
+ N_X_c_314_n N_X_c_303_n N_X_c_317_n N_X_c_304_n N_X_c_330_n N_X_c_306_n
+ N_X_c_310_n N_X_c_312_n Vss PM_G3_DFFQ1_N3_X
x_PM_G3_DFFQ1_N3_Q N_Q_XI4.X0_D N_Q_XI5.X0_D N_Q_c_349_n Q Vss PM_G3_DFFQ1_N3_Q
cc_1 N_VSS_XI1.X0_PGS N_CK_XI13.X0_PGS 0.00316278f
cc_2 N_VSS_XI13.X0_PGD N_CK_XI13.X0_PGS 0.00164185f
cc_3 N_VSS_c_3_p N_CK_XI13.X0_PGS 8.34822e-19
cc_4 N_VSS_c_4_p N_CK_XI13.X0_PGS 4.02129e-19
cc_5 N_VSS_XI1.X0_PGD N_CK_c_106_n 4.20343e-19
cc_6 N_VSS_XI1.X0_PGS N_CK_c_107_n 4.31283e-19
cc_7 N_VSS_c_7_p CK 5.33707e-19
cc_8 N_VSS_XI1.X0_PGD N_VDD_XI0.X0_PGD 0.00196344f
cc_9 N_VSS_XI5.X0_PGD N_VDD_XI4.X0_PGD 0.00221489f
cc_10 N_VSS_XI13.X0_PGD N_VDD_XI12.X0_PGD 0.00211593f
cc_11 N_VSS_c_11_p N_VDD_c_138_n 0.00196344f
cc_12 N_VSS_c_12_p N_VDD_c_139_n 0.00221489f
cc_13 N_VSS_c_13_p N_VDD_c_140_n 0.00211593f
cc_14 N_VSS_c_14_p N_VDD_c_141_n 9.5668e-19
cc_15 N_VSS_c_15_p N_VDD_c_141_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_141_n 0.00423852f
cc_17 N_VSS_c_17_p N_VDD_c_141_n 0.00186049f
cc_18 N_VSS_c_15_p N_VDD_c_145_n 3.48826e-19
cc_19 N_VSS_c_7_p N_VDD_c_145_n 0.00955259f
cc_20 N_VSS_c_20_p N_VDD_c_147_n 0.00105775f
cc_21 N_VSS_c_21_p N_VDD_c_148_n 0.00233232f
cc_22 N_VSS_c_4_p N_VDD_c_148_n 9.47758e-19
cc_23 N_VSS_c_13_p N_VDD_c_150_n 3.69367e-19
cc_24 N_VSS_c_21_p N_VDD_c_150_n 0.00161703f
cc_25 N_VSS_c_4_p N_VDD_c_150_n 2.24973e-19
cc_26 N_VSS_c_7_p N_VDD_c_150_n 0.00142089f
cc_27 N_VSS_c_27_p N_VDD_c_150_n 0.00431851f
cc_28 N_VSS_c_28_p N_VDD_c_150_n 7.74609e-19
cc_29 N_VSS_c_3_p N_VDD_c_156_n 0.00179097f
cc_30 N_VSS_c_30_p N_VDD_c_156_n 3.92901e-19
cc_31 N_VSS_c_31_p N_VDD_c_156_n 8.83788e-19
cc_32 N_VSS_c_12_p N_VDD_c_159_n 3.71132e-19
cc_33 N_VSS_c_31_p N_VDD_c_159_n 0.00141228f
cc_34 N_VSS_c_34_p N_VDD_c_159_n 0.00114511f
cc_35 N_VSS_c_35_p N_VDD_c_159_n 0.00431473f
cc_36 N_VSS_c_36_p N_VDD_c_159_n 0.00338293f
cc_37 N_VSS_c_37_p N_VDD_c_159_n 7.74609e-19
cc_38 N_VSS_c_35_p N_VDD_c_165_n 0.00147849f
cc_39 N_VSS_c_21_p N_VDD_c_166_n 9.29349e-19
cc_40 N_VSS_c_4_p N_VDD_c_166_n 3.79458e-19
cc_41 N_VSS_c_41_p N_VDD_c_168_n 2.72411e-19
cc_42 N_VSS_c_42_p N_VDD_c_168_n 3.23198e-19
cc_43 N_VSS_c_27_p N_VDD_c_168_n 0.00448754f
cc_44 N_VSS_c_44_p N_VDD_c_171_n 4.01154e-19
cc_45 N_VSS_c_42_p N_VDD_c_172_n 0.00187494f
cc_46 N_VSS_c_46_p N_VDD_c_172_n 0.00427673f
cc_47 N_VSS_c_47_p N_VDD_c_172_n 0.00924147f
cc_48 N_VSS_c_48_p N_VDD_c_172_n 9.16632e-19
cc_49 N_VSS_c_31_p N_VDD_c_176_n 4.35319e-19
cc_50 N_VSS_c_34_p N_VDD_c_176_n 4.7255e-19
cc_51 N_VSS_c_36_p N_VDD_c_176_n 0.00107125f
cc_52 N_VSS_c_47_p N_VDD_c_176_n 0.00412661f
cc_53 N_VSS_c_3_p N_VDD_c_180_n 6.19689e-19
cc_54 N_VSS_c_54_p N_VDD_c_180_n 3.8721e-19
cc_55 N_VSS_c_15_p N_VDD_c_182_n 0.00178973f
cc_56 N_VSS_c_7_p N_VDD_c_182_n 2.411e-19
cc_57 N_VSS_c_7_p N_VDD_c_184_n 0.00122269f
cc_58 N_VSS_c_27_p N_VDD_c_185_n 0.00106206f
cc_59 N_VSS_c_47_p N_VDD_c_186_n 0.00116512f
cc_60 N_VSS_c_3_p N_VDD_c_187_n 3.86162e-19
cc_61 N_VSS_c_54_p N_VDD_c_187_n 6.0892e-19
cc_62 N_VSS_c_3_p N_VDD_c_189_n 5.2607e-19
cc_63 N_VSS_c_31_p N_VDD_c_189_n 3.48267e-19
cc_64 N_VSS_c_34_p N_VDD_c_189_n 6.489e-19
cc_65 N_VSS_c_21_p N_VDD_c_192_n 3.48267e-19
cc_66 N_VSS_c_4_p N_VDD_c_192_n 6.20986e-19
cc_67 N_VSS_c_14_p N_CKN_c_242_n 3.43419e-19
cc_68 N_VSS_c_15_p N_CKN_c_242_n 3.48267e-19
cc_69 N_VSS_c_15_p N_CKN_c_244_n 0.00109746f
cc_70 N_VSS_c_3_p N_CKN_c_244_n 6.97825e-19
cc_71 N_VSS_c_7_p N_CKN_c_244_n 3.92176e-19
cc_72 N_VSS_c_47_p N_CKN_c_244_n 3.27346e-19
cc_73 N_VSS_c_47_p N_CKN_c_248_n 0.00111539f
cc_74 N_VSS_c_3_p N_CKN_c_249_n 0.00232042f
cc_75 N_VSS_c_30_p N_CKN_c_249_n 5.94801e-19
cc_76 N_VSS_c_31_p N_CKN_c_249_n 3.31491e-19
cc_77 N_VSS_c_7_p N_CKN_c_249_n 0.00107666f
cc_78 N_VSS_c_78_p N_CKN_c_249_n 5.98734e-19
cc_79 N_VSS_c_35_p N_CKN_c_249_n 6.19556e-19
cc_80 N_VSS_c_27_p N_CKN_c_249_n 7.49546e-19
cc_81 N_VSS_c_81_p N_D_c_279_n 5.28294e-19
cc_82 N_VSS_XI13.X0_PGD N_D_c_280_n 3.99797e-19
cc_83 N_VSS_c_3_p N_D_c_281_n 6.13924e-19
cc_84 N_VSS_c_54_p N_D_c_281_n 3.48267e-19
cc_85 N_VSS_c_4_p N_D_c_281_n 2.1322e-19
cc_86 N_VSS_c_3_p N_D_c_284_n 3.48267e-19
cc_87 N_VSS_c_21_p N_D_c_284_n 2.1322e-19
cc_88 N_VSS_c_54_p N_D_c_284_n 6.88619e-19
cc_89 N_VSS_XI5.X0_PGD N_X_c_303_n 4.09718e-19
cc_90 N_VSS_c_41_p N_X_c_304_n 3.43419e-19
cc_91 N_VSS_c_42_p N_X_c_304_n 3.48267e-19
cc_92 N_VSS_c_41_p N_X_c_306_n 3.48267e-19
cc_93 N_VSS_c_3_p N_X_c_306_n 4.71026e-19
cc_94 N_VSS_c_42_p N_X_c_306_n 5.71987e-19
cc_95 N_VSS_c_47_p N_X_c_306_n 3.92273e-19
cc_96 N_VSS_c_3_p N_X_c_310_n 0.00157847f
cc_97 N_VSS_c_47_p N_X_c_310_n 2.88807e-19
cc_98 N_VSS_c_3_p N_X_c_312_n 3.48267e-19
cc_99 N_VSS_c_99_p N_Q_c_349_n 3.43419e-19
cc_100 N_VSS_c_30_p N_Q_c_349_n 3.48267e-19
cc_101 N_VSS_c_30_p Q 5.37696e-19
cc_102 N_CK_c_106_n N_VDD_XI0.X0_PGD 4.20343e-19
cc_103 N_CK_XI13.X0_PGS N_VDD_XI12.X0_PGD 2.44781e-19
cc_104 N_CK_c_107_n N_VDD_c_140_n 2.44781e-19
cc_105 N_CK_c_107_n N_VDD_c_197_n 2.19802e-19
cc_106 CK N_VDD_c_141_n 5.04211e-19
cc_107 N_CK_c_114_p N_VDD_c_141_n 5.29229e-19
cc_108 N_CK_c_106_n N_VDD_c_145_n 0.00150929f
cc_109 CK N_VDD_c_145_n 0.00141439f
cc_110 N_CK_c_114_p N_VDD_c_145_n 0.0012022f
cc_111 N_CK_XI13.X0_PGS N_VDD_c_148_n 2.48209e-19
cc_112 N_CK_c_107_n N_VDD_c_148_n 5.56076e-19
cc_113 CK N_VDD_c_148_n 3.85155e-19
cc_114 N_CK_c_114_p N_VDD_c_148_n 2.72301e-19
cc_115 CK N_VDD_c_180_n 2.86209e-19
cc_116 N_CK_c_114_p N_VDD_c_180_n 2.18105e-19
cc_117 N_CK_c_124_p N_VDD_c_187_n 5.26604e-19
cc_118 CK N_VDD_c_187_n 2.1322e-19
cc_119 N_CK_XI13.X0_PGS N_CKN_XI12.X0_PGS 4.11563e-19
cc_120 N_CK_XI13.X0_PGS N_CKN_c_257_n 2.73384e-19
cc_121 N_CK_c_106_n N_CKN_c_242_n 7.69306e-19
cc_122 N_CK_XI13.X0_PGS N_D_XI13.X0_CG 4.28946e-19
cc_123 N_CK_XI13.X0_PGS N_D_XI12.X0_CG 2.59344e-19
cc_124 N_CK_XI13.X0_PGS N_D_c_284_n 0.00300565f
cc_125 N_CK_XI13.X0_PGS N_X_XI5.X0_CG 2.61247e-19
cc_126 N_CK_XI13.X0_PGS N_X_c_314_n 4.55333e-19
cc_127 N_CK_XI13.X0_PGS N_X_c_312_n 0.00630896f
cc_128 N_VDD_c_172_n N_CKN_XI12.X0_PGS 8.30122e-19
cc_129 N_VDD_c_172_n N_CKN_c_257_n 8.21431e-19
cc_130 N_VDD_c_197_n N_CKN_c_242_n 3.43419e-19
cc_131 N_VDD_c_145_n N_CKN_c_242_n 2.72411e-19
cc_132 N_VDD_c_197_n N_CKN_c_244_n 3.48267e-19
cc_133 N_VDD_c_141_n N_CKN_c_244_n 6.86019e-19
cc_134 N_VDD_c_145_n N_CKN_c_244_n 2.91445e-19
cc_135 N_VDD_c_148_n N_CKN_c_244_n 5.37696e-19
cc_136 N_VDD_c_180_n N_CKN_c_244_n 6.42405e-19
cc_137 N_VDD_c_172_n N_CKN_c_248_n 7.71262e-19
cc_138 N_VDD_c_166_n N_CKN_c_249_n 2.24632e-19
cc_139 N_VDD_XI12.X0_PGD N_D_c_280_n 4.09718e-19
cc_140 N_VDD_XI4.X0_PGD N_X_c_303_n 3.98597e-19
cc_141 N_VDD_c_224_p N_X_c_317_n 4.97416e-19
cc_142 N_VDD_c_197_n N_X_c_304_n 3.43419e-19
cc_143 N_VDD_c_148_n N_X_c_304_n 3.48267e-19
cc_144 N_VDD_c_150_n N_X_c_304_n 2.72411e-19
cc_145 N_VDD_c_197_n N_X_c_306_n 3.48267e-19
cc_146 N_VDD_c_148_n N_X_c_306_n 6.94315e-19
cc_147 N_VDD_c_150_n N_X_c_306_n 3.78778e-19
cc_148 N_VDD_c_172_n N_X_c_306_n 0.00131866f
cc_149 N_VDD_c_156_n N_X_c_310_n 2.90053e-19
cc_150 N_VDD_c_172_n N_X_c_310_n 2.02855e-19
cc_151 N_VDD_c_189_n N_X_c_310_n 2.26379e-19
cc_152 N_VDD_c_156_n N_X_c_312_n 2.28697e-19
cc_153 N_VDD_c_236_p N_Q_c_349_n 3.43419e-19
cc_154 N_VDD_c_159_n N_Q_c_349_n 2.74986e-19
cc_155 N_VDD_c_171_n N_Q_c_349_n 3.72199e-19
cc_156 N_VDD_c_236_p Q 3.48267e-19
cc_157 N_VDD_c_159_n Q 3.66281e-19
cc_158 N_VDD_c_171_n Q 7.06537e-19
cc_159 N_CKN_XI12.X0_PGS N_D_XI12.X0_CG 0.00419505f
cc_160 N_CKN_c_249_n N_D_c_281_n 2.01502e-19
cc_161 N_CKN_XI12.X0_PGS N_X_c_303_n 0.00422719f
cc_162 N_CKN_c_257_n N_X_c_330_n 5.71169e-19
cc_163 N_CKN_c_249_n N_X_c_330_n 0.00194262f
cc_164 N_CKN_c_244_n N_X_c_306_n 7.35688e-19
cc_165 N_CKN_c_248_n N_X_c_306_n 8.08281e-19
cc_166 N_CKN_c_249_n N_X_c_306_n 7.34542e-19
cc_167 N_CKN_c_249_n N_X_c_310_n 8.56658e-19
cc_168 N_D_c_280_n N_X_c_303_n 0.00477695f
cc_169 N_D_c_280_n N_X_c_304_n 6.90199e-19
cc_170 N_D_c_280_n N_X_c_330_n 4.21501e-19
cc_171 N_D_c_280_n N_X_c_306_n 3.40033e-19
cc_172 N_D_c_281_n N_X_c_306_n 0.00151909f
cc_173 N_D_c_284_n N_X_c_306_n 0.00104518f
cc_174 N_D_c_281_n N_X_c_310_n 0.00146206f
cc_175 N_D_c_284_n N_X_c_310_n 0.00103457f
cc_176 N_D_c_281_n N_X_c_312_n 4.56568e-19
cc_177 N_D_c_284_n N_X_c_312_n 0.00383269f
cc_178 N_X_c_303_n N_Q_c_349_n 6.90199e-19
cc_179 N_X_c_330_n N_Q_c_349_n 3.5757e-19
cc_180 N_X_c_330_n Q 5.52904e-19
*
.ends
*
*
.subckt DFFQ1_HPNW12 CK D Q VDD VSS
xgate (VSS CK VDD D Q) G3_DFFQ1_N3
.ends
*
* File: G1_INV1_N3.pex.netlist
* Created: Fri Feb 25 16:26:51 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G1_INV1_N3_VDD 2 5 15 23 28 30 34 37 43 Vss
c22 43 Vss 0.00440656f
c23 34 Vss 7.98732e-19
c24 30 Vss 0.00491201f
c25 28 Vss 0.0026398f
c26 26 Vss 0.00168274f
c27 23 Vss 0.00814922f
c28 15 Vss 0.0356247f
c29 14 Vss 0.102427f
c30 5 Vss 0.382574f
r31 34 43 1.16709
r32 32 34 2.41736
r33 31 37 0.326018
r34 30 32 0.652036
r35 30 31 7.46046
r36 26 37 0.326018
r37 26 28 6.4185
r38 23 28 1.16709
r39 17 43 0.0476429
r40 15 17 1.45875
r41 14 18 0.652036
r42 14 17 1.45875
r43 11 15 0.652036
r44 5 18 5.1348
r45 5 11 5.1348
r46 2 23 0.123773
.ends

.subckt PM_G1_INV1_N3_A 2 4 12 24 27 Vss
c6 27 Vss 0.00733896f
c7 24 Vss 1.81646e-19
c8 12 Vss 0.229828f
c9 9 Vss 0.180667f
c10 7 Vss 0.0247918f
c11 4 Vss 0.193588f
r12 24 27 1.16709
r13 15 27 0.0476429
r14 13 15 0.326018
r15 13 15 0.1167
r16 12 16 0.652036
r17 12 15 6.7686
r18 9 27 0.357321
r19 7 15 0.326018
r20 7 9 0.40845
r21 4 16 5.1348
r22 2 9 4.72635
.ends

.subckt PM_G1_INV1_N3_VSS 3 6 14 24 27 32 37 49 50 56 Vss
c23 51 Vss 0.0012698f
c24 50 Vss 6.56512e-19
c25 49 Vss 0.00353949f
c26 37 Vss 0.00390919f
c27 32 Vss 0.00198602f
c28 27 Vss 8.43451e-19
c29 24 Vss 0.0100686f
c30 15 Vss 0.0359156f
c31 14 Vss 0.0994171f
c32 3 Vss 0.381612f
r33 51 56 0.326018
r34 49 56 0.326018
r35 49 50 7.46046
r36 45 50 0.652036
r37 32 51 6.4185
r38 27 37 1.16709
r39 27 45 2.41736
r40 24 32 1.16709
r41 17 37 0.0476429
r42 15 17 1.45875
r43 14 18 0.652036
r44 14 17 1.45875
r45 11 15 0.652036
r46 6 24 0.123773
r47 3 18 5.1348
r48 3 11 5.1348
.ends

.subckt PM_G1_INV1_N3_Z 2 4 13 19 Vss
c11 13 Vss 0.00499164f
c12 4 Vss 0.00143493f
r13 16 19 0.0364688
r14 13 16 1.16709
r15 4 13 0.123773
r16 2 13 0.123773
.ends

.subckt G1_INV1_N3  VDD A VSS Z
*
* Z	Z
* VSS	VSS
* A	A
* VDD	VDD
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_A_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW12
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_VSS_XI5.X0_S TIGFET_HPNW12
*
x_PM_G1_INV1_N3_VDD N_VDD_XI6.X0_S N_VDD_XI5.X0_PGD N_VDD_c_4_p N_VDD_c_17_p
+ N_VDD_c_3_p N_VDD_c_5_p N_VDD_c_8_p VDD N_VDD_c_9_p Vss PM_G1_INV1_N3_VDD
x_PM_G1_INV1_N3_A N_A_XI6.X0_CG N_A_XI5.X0_CG N_A_c_23_n A N_A_c_26_p Vss
+ PM_G1_INV1_N3_A
x_PM_G1_INV1_N3_VSS N_VSS_XI6.X0_PGD N_VSS_XI5.X0_S N_VSS_c_31_n N_VSS_c_48_p
+ N_VSS_c_33_n N_VSS_c_37_n N_VSS_c_39_n N_VSS_c_42_n N_VSS_c_43_n VSS Vss
+ PM_G1_INV1_N3_VSS
x_PM_G1_INV1_N3_Z N_Z_XI6.X0_D N_Z_XI5.X0_D N_Z_c_52_n Z Vss PM_G1_INV1_N3_Z
cc_1 N_VDD_XI5.X0_PGD N_A_c_23_n 4.31283e-19
cc_2 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.00199939f
cc_3 N_VDD_c_3_p N_VSS_XI6.X0_PGD 4.23795e-19
cc_4 N_VDD_c_4_p N_VSS_c_31_n 0.00199939f
cc_5 N_VDD_c_5_p N_VSS_c_31_n 5.08727e-19
cc_6 N_VDD_c_3_p N_VSS_c_33_n 0.00302944f
cc_7 N_VDD_c_5_p N_VSS_c_33_n 0.00141897f
cc_8 N_VDD_c_8_p N_VSS_c_33_n 9.31072e-19
cc_9 N_VDD_c_9_p N_VSS_c_33_n 3.48267e-19
cc_10 N_VDD_c_3_p N_VSS_c_37_n 7.58061e-19
cc_11 N_VDD_c_8_p N_VSS_c_37_n 0.00105766f
cc_12 N_VDD_c_3_p N_VSS_c_39_n 9.55109e-19
cc_13 N_VDD_c_5_p N_VSS_c_39_n 0.00103739f
cc_14 N_VDD_c_9_p N_VSS_c_39_n 6.46219e-19
cc_15 N_VDD_c_5_p N_VSS_c_42_n 0.0059288f
cc_16 N_VDD_c_5_p N_VSS_c_43_n 0.00172731f
cc_17 N_VDD_c_17_p N_Z_c_52_n 3.43419e-19
cc_18 N_VDD_c_3_p N_Z_c_52_n 3.48267e-19
cc_19 N_VDD_c_5_p N_Z_c_52_n 2.60012e-19
cc_20 N_VDD_c_17_p Z 3.48267e-19
cc_21 N_VDD_c_3_p Z 7.09569e-19
cc_22 N_VDD_c_5_p Z 3.45966e-19
cc_23 N_A_c_23_n N_VSS_XI6.X0_PGD 4.31283e-19
cc_24 A N_VSS_c_33_n 3.42414e-19
cc_25 N_A_c_26_p N_VSS_c_33_n 2.30774e-19
cc_26 A N_VSS_c_39_n 2.30774e-19
cc_27 N_A_c_23_n N_Z_c_52_n 7.69306e-19
cc_28 N_VSS_c_48_p N_Z_c_52_n 3.43419e-19
cc_29 N_VSS_c_37_n N_Z_c_52_n 3.48267e-19
cc_30 N_VSS_c_37_n Z 8.23589e-19
cc_31 N_VSS_c_42_n Z 2.18525e-19
*
.ends
*
*
.subckt INV1_HPNW12 A Y VDD VSS
xgate (VDD A VSS Y) G1_INV1_N3
.ends
*
* File: G3_LATQ1_N3.pex.netlist
* Created: Tue Apr  5 12:00:00 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_LATQ1_N3_VDD 2 4 6 8 10 12 14 16 31 42 48 58 63 66 68 69 70 71 72
+ 75 77 81 85 90 92 98 103 Vss
c82 103 Vss 0.00476181f
c83 98 Vss 0.00486653f
c84 90 Vss 2.39889e-19
c85 85 Vss 0.00253232f
c86 83 Vss 0.0017055f
c87 81 Vss 0.00108379f
c88 77 Vss 0.0043713f
c89 75 Vss 8.9379e-19
c90 72 Vss 8.65746e-19
c91 71 Vss 0.00223415f
c92 70 Vss 8.64769e-19
c93 69 Vss 0.00576876f
c94 68 Vss 0.0113641f
c95 66 Vss 0.00582672f
c96 63 Vss 0.00607435f
c97 58 Vss 0.00819566f
c98 53 Vss 0.0307825f
c99 48 Vss 0.230506f
c100 44 Vss 1.68267e-19
c101 42 Vss 0.0357228f
c102 41 Vss 0.0656875f
c103 32 Vss 0.0359366f
c104 31 Vss 0.101312f
c105 16 Vss 0.00143493f
c106 14 Vss 0.191707f
c107 10 Vss 0.191287f
c108 8 Vss 0.189707f
c109 6 Vss 0.190072f
c110 4 Vss 0.189718f
r111 83 92 0.326018
r112 83 85 6.16843
r113 81 103 1.16709
r114 79 81 2.16729
r115 78 90 0.494161
r116 77 92 0.326018
r117 77 78 7.46046
r118 75 98 1.16709
r119 73 90 0.128424
r120 73 75 2.16729
r121 71 90 0.494161
r122 71 72 4.37625
r123 69 79 0.652036
r124 69 70 10.1279
r125 68 72 0.652036
r126 67 68 18.2969
r127 66 89 2.334
r128 66 67 0.14525
r129 65 70 0.652036
r130 65 66 5.54325
r131 63 85 1.16709
r132 58 89 1.16709
r133 49 53 0.494161
r134 48 50 0.652036
r135 48 49 6.8853
r136 45 53 0.128424
r137 44 103 0.0476429
r138 42 44 1.45875
r139 41 53 0.494161
r140 41 44 1.45875
r141 38 42 0.652036
r142 34 98 0.0476429
r143 32 34 1.45875
r144 31 35 0.652036
r145 31 34 1.45875
r146 28 32 0.652036
r147 16 63 0.123773
r148 14 50 5.1348
r149 12 63 0.123773
r150 10 45 5.1348
r151 8 38 5.1348
r152 6 28 5.1348
r153 4 35 5.1348
r154 2 58 0.123773
.ends

.subckt PM_G3_LATQ1_N3_VSS 2 4 6 8 10 12 14 16 31 32 34 42 48 58 63 66 71 76 81
+ 90 95 104 106 107 108 113 114 119 129 130 132 Vss
c74 130 Vss 3.75522e-19
c75 129 Vss 4.28045e-19
c76 125 Vss 0.00128551f
c77 119 Vss 0.00327372f
c78 114 Vss 8.25631e-19
c79 113 Vss 0.00434469f
c80 108 Vss 8.30816e-19
c81 107 Vss 0.00172205f
c82 106 Vss 0.00206535f
c83 104 Vss 0.00621153f
c84 95 Vss 0.00443295f
c85 90 Vss 0.0041985f
c86 81 Vss 0.00249073f
c87 76 Vss 9.5519e-19
c88 71 Vss 6.07136e-19
c89 66 Vss 0.0013933f
c90 63 Vss 0.0060193f
c91 58 Vss 0.00814768f
c92 53 Vss 0.0307825f
c93 48 Vss 0.231473f
c94 42 Vss 0.0348714f
c95 41 Vss 0.0647879f
c96 34 Vss 8.95828e-20
c97 32 Vss 0.0350852f
c98 31 Vss 0.0994129f
c99 16 Vss 0.191895f
c100 14 Vss 0.00143493f
c101 12 Vss 0.19162f
c102 10 Vss 0.189706f
c103 4 Vss 0.190073f
c104 2 Vss 0.18972f
r105 125 132 0.326018
r106 120 130 0.494161
r107 119 132 0.326018
r108 119 120 7.46046
r109 115 130 0.128424
r110 113 121 0.652036
r111 113 114 10.1279
r112 109 129 0.0828784
r113 107 130 0.494161
r114 107 108 4.37625
r115 106 114 0.652036
r116 105 129 0.551426
r117 105 106 5.50157
r118 104 129 0.551426
r119 103 108 0.652036
r120 103 104 18.3386
r121 81 125 6.16843
r122 76 95 1.16709
r123 76 121 2.16729
r124 71 90 1.16709
r125 71 115 2.16729
r126 66 109 1.82344
r127 63 81 1.16709
r128 58 66 1.16709
r129 49 53 0.494161
r130 48 50 0.652036
r131 48 49 6.8853
r132 45 53 0.128424
r133 44 95 0.0476429
r134 42 44 1.45875
r135 41 53 0.494161
r136 41 44 1.45875
r137 38 42 0.652036
r138 34 90 0.0476429
r139 32 34 1.45875
r140 31 35 0.652036
r141 31 34 1.45875
r142 28 32 0.652036
r143 16 50 5.1348
r144 14 63 0.123773
r145 12 45 5.1348
r146 10 38 5.1348
r147 8 63 0.123773
r148 6 58 0.123773
r149 4 28 5.1348
r150 2 35 5.1348
.ends

.subckt PM_G3_LATQ1_N3_G 2 4 6 14 15 22 31 37 Vss
c24 37 Vss 0.00266632f
c25 31 Vss 6.62558e-19
c26 29 Vss 0.0295325f
c27 22 Vss 0.152777f
c28 15 Vss 0.179526f
c29 14 Vss 2.0264e-19
c30 10 Vss 0.0247918f
c31 6 Vss 0.192371f
c32 4 Vss 0.193138f
c33 2 Vss 0.180487f
r34 34 37 1.16709
r35 31 34 0.0833571
r36 23 29 0.494161
r37 22 24 0.652036
r38 22 23 4.84305
r39 19 29 0.128424
r40 18 37 0.0476429
r41 16 18 0.326018
r42 16 18 0.1167
r43 15 29 0.494161
r44 15 18 6.7686
r45 14 37 0.357321
r46 10 18 0.326018
r47 10 14 0.40845
r48 6 24 5.1348
r49 4 19 5.1348
r50 2 14 4.72635
.ends

.subckt PM_G3_LATQ1_N3_QN 2 4 6 8 20 23 33 37 40 45 48 53 69 Vss
c43 69 Vss 4.86032e-19
c44 53 Vss 0.00238508f
c45 48 Vss 0.00856405f
c46 45 Vss 0.00518251f
c47 40 Vss 0.00103774f
c48 37 Vss 0.0113402f
c49 33 Vss 0.0113402f
c50 23 Vss 2.25442e-19
c51 20 Vss 0.214677f
c52 17 Vss 0.180502f
c53 15 Vss 0.0247918f
c54 4 Vss 0.191818f
r55 65 69 0.652036
r56 48 69 13.7956
r57 48 50 6.4185
r58 45 48 6.4185
r59 40 53 1.16709
r60 40 65 1.83386
r61 37 50 1.16709
r62 33 45 1.16709
r63 23 53 0.0476429
r64 21 23 0.326018
r65 21 23 0.1167
r66 20 24 0.652036
r67 20 23 6.7686
r68 17 53 0.357321
r69 15 23 0.326018
r70 15 17 0.40845
r71 8 37 0.123773
r72 6 33 0.123773
r73 4 24 5.1348
r74 2 17 4.72635
.ends

.subckt PM_G3_LATQ1_N3_GN 2 4 6 12 23 27 29 30 32 39 Vss
c39 39 Vss 0.00500045f
c40 32 Vss 6.08951e-19
c41 30 Vss 6.08791e-19
c42 29 Vss 0.00111596f
c43 27 Vss 0.00109183f
c44 23 Vss 0.00525048f
c45 14 Vss 1.82689e-19
c46 12 Vss 0.163012f
c47 6 Vss 0.285833f
c48 4 Vss 0.00143493f
r49 32 39 1.16709
r50 29 32 0.531835
r51 29 30 1.70882
r52 25 30 0.652036
r53 25 27 5.835
r54 23 27 1.16709
r55 14 39 0.197068
r56 12 16 0.652036
r57 12 14 4.668
r58 6 16 8.4024
r59 4 23 0.123773
r60 2 23 0.123773
.ends

.subckt PM_G3_LATQ1_N3_Q 2 4 13 18 Vss
c12 18 Vss 3.21524e-19
c13 13 Vss 0.00454527f
c14 4 Vss 0.00143493f
r15 13 18 1.16709
r16 4 13 0.123773
r17 2 13 0.123773
.ends

.subckt PM_G3_LATQ1_N3_D 2 4 10 14 Vss
c14 14 Vss 4.85129e-19
c15 10 Vss 1.35847e-19
c16 2 Vss 0.58413f
r17 14 17 0.0416786
r18 10 17 1.16709
r19 4 10 8.9859
r20 2 10 8.9859
.ends

.subckt G3_LATQ1_N3  VDD VSS G Q D
*
* D	D
* Q	Q
* G	G
* VSS	VSS
* VDD	VDD
XI3.X0 N_GN_XI3.X0_D N_VSS_XI3.X0_PGD N_G_XI3.X0_CG N_VSS_XI3.X0_PGS
+ N_VDD_XI3.X0_S TIGFET_HPNW12
XI0.X0 N_Q_XI0.X0_D N_VDD_XI0.X0_PGD N_QN_XI0.X0_CG N_VDD_XI0.X0_PGS
+ N_VSS_XI0.X0_S TIGFET_HPNW12
XI1.X0 N_GN_XI1.X0_D N_VDD_XI1.X0_PGD N_G_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW12
XI4.X0 N_Q_XI4.X0_D N_VSS_XI4.X0_PGD N_QN_XI4.X0_CG N_VSS_XI4.X0_PGS
+ N_VDD_XI4.X0_S TIGFET_HPNW12
XI2.X0 N_QN_XI2.X0_D N_VDD_XI2.X0_PGD N_D_XI2.X0_CG N_G_XI2.X0_PGS
+ N_VSS_XI2.X0_S TIGFET_HPNW12
XI5.X0 N_QN_XI5.X0_D N_VSS_XI5.X0_PGD N_D_XI5.X0_CG N_GN_XI5.X0_PGS
+ N_VDD_XI5.X0_S TIGFET_HPNW12
*
x_PM_G3_LATQ1_N3_VDD N_VDD_XI3.X0_S N_VDD_XI0.X0_PGD N_VDD_XI0.X0_PGS
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI4.X0_S N_VDD_XI2.X0_PGD
+ N_VDD_XI5.X0_S N_VDD_c_9_p N_VDD_c_5_p N_VDD_c_14_p N_VDD_c_69_p N_VDD_c_11_p
+ N_VDD_c_7_p N_VDD_c_13_p N_VDD_c_6_p N_VDD_c_41_p N_VDD_c_18_p N_VDD_c_45_p
+ N_VDD_c_23_p N_VDD_c_10_p N_VDD_c_21_p N_VDD_c_12_p N_VDD_c_44_p VDD
+ N_VDD_c_26_p N_VDD_c_22_p Vss PM_G3_LATQ1_N3_VDD
x_PM_G3_LATQ1_N3_VSS N_VSS_XI3.X0_PGD N_VSS_XI3.X0_PGS N_VSS_XI0.X0_S
+ N_VSS_XI1.X0_S N_VSS_XI4.X0_PGD N_VSS_XI4.X0_PGS N_VSS_XI2.X0_S
+ N_VSS_XI5.X0_PGD N_VSS_c_87_n N_VSS_c_89_n N_VSS_c_131_p N_VSS_c_91_n
+ N_VSS_c_93_n N_VSS_c_95_n N_VSS_c_96_n N_VSS_c_98_n N_VSS_c_101_n
+ N_VSS_c_105_n N_VSS_c_109_n N_VSS_c_111_n N_VSS_c_115_n N_VSS_c_119_n
+ N_VSS_c_121_n N_VSS_c_122_n N_VSS_c_123_n N_VSS_c_124_n N_VSS_c_127_n
+ N_VSS_c_128_n N_VSS_c_129_n N_VSS_c_130_n VSS Vss PM_G3_LATQ1_N3_VSS
x_PM_G3_LATQ1_N3_G N_G_XI3.X0_CG N_G_XI1.X0_CG N_G_XI2.X0_PGS N_G_c_162_n
+ N_G_c_158_n N_G_c_159_n G N_G_c_161_n Vss PM_G3_LATQ1_N3_G
x_PM_G3_LATQ1_N3_QN N_QN_XI0.X0_CG N_QN_XI4.X0_CG N_QN_XI2.X0_D N_QN_XI5.X0_D
+ N_QN_c_181_n N_QN_c_182_n N_QN_c_196_n N_QN_c_183_n N_QN_c_185_n N_QN_c_187_n
+ N_QN_c_189_n N_QN_c_192_n N_QN_c_194_n Vss PM_G3_LATQ1_N3_QN
x_PM_G3_LATQ1_N3_GN N_GN_XI3.X0_D N_GN_XI1.X0_D N_GN_XI5.X0_PGS N_GN_c_224_n
+ N_GN_c_225_n N_GN_c_228_n N_GN_c_244_n N_GN_c_250_n N_GN_c_252_n N_GN_c_245_n
+ Vss PM_G3_LATQ1_N3_GN
x_PM_G3_LATQ1_N3_Q N_Q_XI0.X0_D N_Q_XI4.X0_D N_Q_c_263_n Q Vss PM_G3_LATQ1_N3_Q
x_PM_G3_LATQ1_N3_D N_D_XI2.X0_CG N_D_XI5.X0_CG N_D_c_280_n D Vss
+ PM_G3_LATQ1_N3_D
cc_1 N_VDD_XI1.X0_PGD N_VSS_XI3.X0_PGD 0.00203852f
cc_2 N_VDD_XI0.X0_PGS N_VSS_XI3.X0_PGS 2.44446e-19
cc_3 N_VDD_XI0.X0_PGD N_VSS_XI4.X0_PGD 0.00203076f
cc_4 N_VDD_XI2.X0_PGD N_VSS_XI5.X0_PGD 2.44446e-19
cc_5 N_VDD_c_5_p N_VSS_c_87_n 0.00203852f
cc_6 N_VDD_c_6_p N_VSS_c_87_n 3.89167e-19
cc_7 N_VDD_c_7_p N_VSS_c_89_n 3.80615e-19
cc_8 N_VDD_c_6_p N_VSS_c_89_n 3.89167e-19
cc_9 N_VDD_c_9_p N_VSS_c_91_n 0.00203076f
cc_10 N_VDD_c_10_p N_VSS_c_91_n 3.00073e-19
cc_11 N_VDD_c_11_p N_VSS_c_93_n 2.19802e-19
cc_12 N_VDD_c_12_p N_VSS_c_93_n 8.58125e-19
cc_13 N_VDD_c_13_p N_VSS_c_95_n 9.5668e-19
cc_14 N_VDD_c_14_p N_VSS_c_96_n 2.19802e-19
cc_15 N_VDD_c_11_p N_VSS_c_96_n 2.80254e-19
cc_16 N_VDD_c_7_p N_VSS_c_98_n 4.06916e-19
cc_17 N_VDD_c_13_p N_VSS_c_98_n 0.00165395f
cc_18 N_VDD_c_18_p N_VSS_c_98_n 3.5277e-19
cc_19 N_VDD_c_7_p N_VSS_c_101_n 9.31121e-19
cc_20 N_VDD_c_6_p N_VSS_c_101_n 0.00161703f
cc_21 N_VDD_c_21_p N_VSS_c_101_n 7.09654e-19
cc_22 N_VDD_c_22_p N_VSS_c_101_n 3.48267e-19
cc_23 N_VDD_c_23_p N_VSS_c_105_n 9.52068e-19
cc_24 N_VDD_c_10_p N_VSS_c_105_n 0.00141228f
cc_25 N_VDD_c_12_p N_VSS_c_105_n 0.00257912f
cc_26 N_VDD_c_26_p N_VSS_c_105_n 3.48267e-19
cc_27 N_VDD_c_7_p N_VSS_c_109_n 3.32876e-19
cc_28 N_VDD_c_21_p N_VSS_c_109_n 8.43845e-19
cc_29 N_VDD_c_7_p N_VSS_c_111_n 4.24454e-19
cc_30 N_VDD_c_6_p N_VSS_c_111_n 2.26455e-19
cc_31 N_VDD_c_21_p N_VSS_c_111_n 3.84769e-19
cc_32 N_VDD_c_22_p N_VSS_c_111_n 6.489e-19
cc_33 N_VDD_c_23_p N_VSS_c_115_n 3.82294e-19
cc_34 N_VDD_c_10_p N_VSS_c_115_n 0.00114511f
cc_35 N_VDD_c_12_p N_VSS_c_115_n 9.55109e-19
cc_36 N_VDD_c_26_p N_VSS_c_115_n 6.46219e-19
cc_37 N_VDD_c_7_p N_VSS_c_119_n 0.00540208f
cc_38 N_VDD_c_13_p N_VSS_c_119_n 0.00786235f
cc_39 N_VDD_c_13_p N_VSS_c_121_n 0.00445899f
cc_40 N_VDD_c_6_p N_VSS_c_122_n 0.00348718f
cc_41 N_VDD_c_41_p N_VSS_c_123_n 0.00106807f
cc_42 N_VDD_c_18_p N_VSS_c_124_n 0.00356332f
cc_43 N_VDD_c_10_p N_VSS_c_124_n 0.00600653f
cc_44 N_VDD_c_44_p N_VSS_c_124_n 0.00103147f
cc_45 N_VDD_c_45_p N_VSS_c_127_n 0.00106428f
cc_46 N_VDD_c_6_p N_VSS_c_128_n 0.00586992f
cc_47 N_VDD_c_13_p N_VSS_c_129_n 9.16632e-19
cc_48 N_VDD_c_6_p N_VSS_c_130_n 7.74609e-19
cc_49 N_VDD_c_14_p N_G_XI2.X0_PGS 0.00172513f
cc_50 N_VDD_XI1.X0_PGD N_G_c_158_n 3.99191e-19
cc_51 N_VDD_XI1.X0_PGS N_G_c_159_n 4.09718e-19
cc_52 N_VDD_c_13_p G 5.04211e-19
cc_53 N_VDD_c_13_p N_G_c_161_n 5.56409e-19
cc_54 N_VDD_XI0.X0_PGD N_QN_c_181_n 4.09718e-19
cc_55 N_VDD_c_26_p N_QN_c_182_n 6.34963e-19
cc_56 N_VDD_c_11_p N_QN_c_183_n 3.43419e-19
cc_57 N_VDD_c_12_p N_QN_c_183_n 3.48267e-19
cc_58 N_VDD_c_13_p N_QN_c_185_n 4.49462e-19
cc_59 N_VDD_c_26_p N_QN_c_185_n 2.10618e-19
cc_60 N_VDD_c_11_p N_QN_c_187_n 3.48267e-19
cc_61 N_VDD_c_12_p N_QN_c_187_n 9.04108e-19
cc_62 N_VDD_c_6_p N_QN_c_189_n 3.28643e-19
cc_63 N_VDD_c_10_p N_QN_c_189_n 2.94643e-19
cc_64 N_VDD_c_12_p N_QN_c_189_n 3.47038e-19
cc_65 N_VDD_c_13_p N_QN_c_192_n 2.92308e-19
cc_66 N_VDD_c_23_p N_QN_c_192_n 2.28697e-19
cc_67 N_VDD_c_13_p N_QN_c_194_n 3.90734e-19
cc_68 N_VDD_c_11_p N_GN_c_224_n 3.11705e-19
cc_69 N_VDD_c_69_p N_GN_c_225_n 3.43419e-19
cc_70 N_VDD_c_7_p N_GN_c_225_n 3.72199e-19
cc_71 N_VDD_c_6_p N_GN_c_225_n 2.74986e-19
cc_72 N_VDD_c_69_p N_GN_c_228_n 3.48267e-19
cc_73 N_VDD_c_7_p N_GN_c_228_n 7.94301e-19
cc_74 N_VDD_c_13_p N_GN_c_228_n 0.00122181f
cc_75 N_VDD_c_6_p N_GN_c_228_n 3.82604e-19
cc_76 N_VDD_c_11_p N_Q_c_263_n 3.43419e-19
cc_77 N_VDD_c_10_p N_Q_c_263_n 2.74986e-19
cc_78 N_VDD_c_12_p N_Q_c_263_n 3.48267e-19
cc_79 N_VDD_c_11_p Q 3.48267e-19
cc_80 N_VDD_c_10_p Q 3.66281e-19
cc_81 N_VDD_c_12_p Q 7.09569e-19
cc_82 N_VDD_c_14_p N_D_XI2.X0_CG 4.32953e-19
cc_83 N_VSS_c_131_p N_G_c_162_n 5.35095e-19
cc_84 N_VSS_XI3.X0_PGD N_G_c_158_n 4.09718e-19
cc_85 N_VSS_c_111_n G 2.15082e-19
cc_86 N_VSS_c_119_n G 2.86445e-19
cc_87 N_VSS_c_101_n N_G_c_161_n 2.15082e-19
cc_88 N_VSS_XI4.X0_PGD N_QN_c_181_n 3.99191e-19
cc_89 N_VSS_c_96_n N_QN_c_196_n 3.43419e-19
cc_90 N_VSS_c_109_n N_QN_c_196_n 3.48267e-19
cc_91 N_VSS_c_96_n N_QN_c_187_n 3.48267e-19
cc_92 N_VSS_c_109_n N_QN_c_187_n 8.62542e-19
cc_93 N_VSS_c_109_n N_QN_c_189_n 5.58212e-19
cc_94 N_VSS_c_124_n N_QN_c_189_n 4.58442e-19
cc_95 N_VSS_c_128_n N_QN_c_189_n 6.13056e-19
cc_96 N_VSS_c_101_n N_QN_c_194_n 3.59967e-19
cc_97 N_VSS_c_119_n N_QN_c_194_n 0.00182171f
cc_98 N_VSS_c_93_n N_GN_XI5.X0_PGS 0.00172853f
cc_99 N_VSS_XI4.X0_PGS N_GN_c_224_n 6.66551e-19
cc_100 N_VSS_c_96_n N_GN_c_225_n 3.43419e-19
cc_101 N_VSS_c_109_n N_GN_c_225_n 3.48267e-19
cc_102 N_VSS_c_96_n N_GN_c_228_n 3.48267e-19
cc_103 N_VSS_c_109_n N_GN_c_228_n 4.99861e-19
cc_104 N_VSS_c_119_n N_GN_c_228_n 7.12611e-19
cc_105 N_VSS_c_95_n N_Q_c_263_n 3.43419e-19
cc_106 N_VSS_c_98_n N_Q_c_263_n 3.48267e-19
cc_107 N_VSS_c_98_n Q 8.15956e-19
cc_108 N_VSS_c_93_n N_D_XI2.X0_CG 4.32953e-19
cc_109 N_G_c_158_n N_QN_c_181_n 0.00400131f
cc_110 G N_QN_c_185_n 4.48861e-19
cc_111 N_G_c_161_n N_QN_c_185_n 4.54925e-19
cc_112 G N_QN_c_192_n 4.56568e-19
cc_113 N_G_c_161_n N_QN_c_192_n 0.00268575f
cc_114 N_G_c_159_n N_GN_c_224_n 0.00878732f
cc_115 N_G_c_158_n N_GN_c_225_n 6.90199e-19
cc_116 N_G_c_158_n N_GN_c_228_n 3.82175e-19
cc_117 G N_GN_c_228_n 0.00151253f
cc_118 N_G_c_161_n N_GN_c_228_n 9.72448e-19
cc_119 N_G_c_158_n N_GN_c_244_n 4.1347e-19
cc_120 N_G_c_158_n N_GN_c_245_n 0.00397074f
cc_121 N_G_c_161_n N_GN_c_245_n 2.41671e-19
cc_122 N_G_XI2.X0_PGS N_D_XI2.X0_CG 0.00435077f
cc_123 N_QN_c_181_n N_GN_XI5.X0_PGS 0.00196434f
cc_124 N_QN_c_187_n N_GN_c_228_n 0.00124016f
cc_125 N_QN_c_189_n N_GN_c_244_n 0.00100851f
cc_126 N_QN_c_181_n N_GN_c_250_n 4.04137e-19
cc_127 N_QN_c_189_n N_GN_c_250_n 0.00133182f
cc_128 N_QN_c_189_n N_GN_c_252_n 0.00102929f
cc_129 N_QN_c_181_n N_GN_c_245_n 0.00341994f
cc_130 N_QN_c_192_n N_GN_c_245_n 2.75519e-19
cc_131 N_QN_c_181_n N_Q_c_263_n 6.90199e-19
cc_132 N_QN_c_181_n N_D_XI2.X0_CG 3.26559e-19
cc_133 N_QN_c_187_n N_D_XI2.X0_CG 0.0010503f
cc_134 N_QN_c_187_n N_D_c_280_n 0.00130556f
cc_135 N_QN_c_187_n D 0.00141415f
cc_136 N_QN_c_189_n D 0.00146947f
cc_137 N_GN_c_250_n N_Q_c_263_n 3.29741e-19
cc_138 N_GN_c_250_n Q 3.9897e-19
cc_139 N_GN_XI5.X0_PGS N_D_XI2.X0_CG 0.0048787f
cc_140 N_GN_c_224_n N_D_c_280_n 0.00333193f
cc_141 N_GN_c_252_n N_D_c_280_n 3.73302e-19
cc_142 N_GN_c_245_n N_D_c_280_n 8.5422e-19
cc_143 N_GN_c_252_n D 2.85187e-19
cc_144 N_GN_c_245_n D 3.48267e-19
*
.ends
*
*
.subckt LATQ1_HPNW12 D G Q VDD VSS
xgate (VDD VSS G Q D) G3_LATQ1_N3
.ends
*
* File: G4_MAJ3_N3.pex.netlist
* Created: Fri Mar  4 11:51:04 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MAJ3_N3_VDD 2 4 7 11 27 28 30 31 32 44 48 52 54 56 57 58 61 65 67
+ 69 70 73 77 79 80 90 95 Vss
c76 95 Vss 0.00472824f
c77 90 Vss 0.00466016f
c78 80 Vss 4.52364e-19
c79 79 Vss 4.28405e-19
c80 77 Vss 4.68316e-19
c81 73 Vss 0.00105057f
c82 70 Vss 8.64769e-19
c83 69 Vss 0.00576436f
c84 67 Vss 0.00145931f
c85 61 Vss 0.00146297f
c86 58 Vss 8.64769e-19
c87 57 Vss 0.00590519f
c88 56 Vss 0.0027558f
c89 54 Vss 0.0069447f
c90 52 Vss 0.00282697f
c91 48 Vss 0.00810125f
c92 44 Vss 0.0099068f
c93 32 Vss 0.0356247f
c94 31 Vss 0.10084f
c95 28 Vss 0.0356247f
c96 27 Vss 0.100978f
c97 11 Vss 0.376343f
c98 7 Vss 0.374237f
r99 77 95 1.16709
r100 75 77 2.16729
r101 73 90 1.16709
r102 71 73 2.16729
r103 69 75 0.652036
r104 69 70 10.1279
r105 65 67 1.167
r106 63 80 0.0828784
r107 63 65 0.656438
r108 59 79 0.0828784
r109 59 61 1.82344
r110 57 71 0.652036
r111 57 58 10.1279
r112 56 70 0.652036
r113 55 80 0.551426
r114 55 56 5.50157
r115 54 80 0.551426
r116 53 79 0.551426
r117 53 54 11.5033
r118 52 79 0.551426
r119 51 58 0.652036
r120 51 52 5.50157
r121 48 67 1.16709
r122 44 61 1.16709
r123 34 95 0.0476429
r124 32 34 1.45875
r125 31 38 0.652036
r126 31 34 1.45875
r127 30 90 0.0476429
r128 28 30 1.45875
r129 27 35 0.652036
r130 27 30 1.45875
r131 24 32 0.652036
r132 21 28 0.652036
r133 11 38 5.1348
r134 11 24 5.1348
r135 7 35 5.1348
r136 7 21 5.1348
r137 4 48 0.123773
r138 2 44 0.123773
.ends

.subckt PM_G4_MAJ3_N3_VSS 3 7 10 12 27 28 31 32 45 49 52 57 62 67 70 73 78 91 92
+ 93 94 95 104 114 115 117 Vss
c81 115 Vss 3.75522e-19
c82 114 Vss 3.75522e-19
c83 110 Vss 0.00128551f
c84 104 Vss 0.00368719f
c85 95 Vss 8.30816e-19
c86 94 Vss 0.00157211f
c87 93 Vss 8.30816e-19
c88 92 Vss 0.00157211f
c89 91 Vss 0.00860014f
c90 78 Vss 0.00407667f
c91 73 Vss 0.00419321f
c92 70 Vss 0.00352694f
c93 67 Vss 0.00278012f
c94 62 Vss 0.00185852f
c95 57 Vss 0.00149825f
c96 52 Vss 0.00105861f
c97 49 Vss 0.00997263f
c98 45 Vss 0.00798745f
c99 32 Vss 0.0350852f
c100 31 Vss 0.0994129f
c101 28 Vss 0.0350852f
c102 27 Vss 0.0994129f
c103 7 Vss 0.377882f
c104 3 Vss 0.379585f
r105 110 117 0.326018
r106 106 115 0.494161
r107 105 114 0.494161
r108 104 117 0.326018
r109 104 105 7.46046
r110 100 115 0.128424
r111 96 114 0.128424
r112 94 115 0.494161
r113 94 95 4.37625
r114 92 114 0.494161
r115 92 93 4.37625
r116 91 95 0.652036
r117 90 93 0.652036
r118 90 91 25.1739
r119 70 106 8.04396
r120 67 70 6.75193
r121 62 110 6.16843
r122 57 78 1.16709
r123 57 100 2.16729
r124 52 73 1.16709
r125 52 96 2.16729
r126 49 67 1.16709
r127 45 62 1.16709
r128 34 78 0.0476429
r129 32 34 1.45875
r130 31 38 0.652036
r131 31 34 1.45875
r132 30 73 0.0476429
r133 28 30 1.45875
r134 27 35 0.652036
r135 27 30 1.45875
r136 24 32 0.652036
r137 21 28 0.652036
r138 12 49 0.123773
r139 10 45 0.123773
r140 7 38 5.1348
r141 7 24 5.1348
r142 3 35 5.1348
r143 3 21 5.1348
.ends

.subckt PM_G4_MAJ3_N3_A 2 4 6 8 11 15 32 53 57 62 67 69 72 74 76 79 81 87 89 97
+ 100 109 Vss
c72 109 Vss 0.00544007f
c73 100 Vss 0.00497933f
c74 97 Vss 1.8079e-19
c75 94 Vss 7.63366e-19
c76 89 Vss 8.03875e-19
c77 87 Vss 8.73696e-19
c78 83 Vss 0.0024194f
c79 81 Vss 0.00445355f
c80 79 Vss 6.95023e-19
c81 76 Vss 0.00110877f
c82 75 Vss 0.00146569f
c83 74 Vss 0.00592189f
c84 69 Vss 0.00755424f
c85 67 Vss 0.0082356f
c86 62 Vss 0.00963114f
c87 57 Vss 0.135088f
c88 53 Vss 0.127963f
c89 32 Vss 0.217507f
c90 29 Vss 0.180502f
c91 27 Vss 0.0247918f
c92 11 Vss 1.44228f
c93 4 Vss 0.193588f
r94 109 112 0.1
r95 97 109 1.16709
r96 92 100 1.16709
r97 89 92 1.08364
r98 85 87 3.501
r99 84 97 0.0685365
r100 83 85 0.652036
r101 83 84 1.70882
r102 82 94 0.494161
r103 81 97 0.0685365
r104 81 82 7.46046
r105 77 94 0.128424
r106 77 79 3.501
r107 75 94 0.494161
r108 75 76 1.83386
r109 73 76 0.652036
r110 73 74 10.6697
r111 70 89 0.0685365
r112 70 72 1.41707
r113 69 74 0.652036
r114 69 72 8.79418
r115 67 87 1.16709
r116 62 79 1.16709
r117 55 57 4.53833
r118 52 112 0.0238214
r119 52 53 2.26917
r120 49 52 2.26917
r121 44 57 0.00605528
r122 43 53 0.00605528
r123 40 55 0.00605528
r124 39 49 0.00605528
r125 35 100 0.0476429
r126 33 35 0.326018
r127 33 35 0.1167
r128 32 36 0.652036
r129 32 35 6.7686
r130 29 100 0.357321
r131 27 35 0.326018
r132 27 29 0.40845
r133 15 44 5.1348
r134 15 40 5.1348
r135 11 15 17.9718
r136 11 43 5.1348
r137 11 15 17.9718
r138 11 39 5.1348
r139 8 67 0.123773
r140 6 62 0.123773
r141 4 36 5.1348
r142 2 29 4.72635
.ends

.subckt PM_G4_MAJ3_N3_BI 2 4 6 8 21 29 32 37 42 52 57 66 72 73 81 Vss
c58 81 Vss 5.35611e-19
c59 73 Vss 2.99365e-19
c60 72 Vss 7.27663e-19
c61 66 Vss 0.00156866f
c62 57 Vss 0.00147096f
c63 52 Vss 0.00166247f
c64 42 Vss 0.00166542f
c65 37 Vss 0.005464f
c66 32 Vss 0.00219142f
c67 29 Vss 0.00514303f
c68 21 Vss 0.166484f
c69 6 Vss 0.166484f
c70 4 Vss 0.00143493f
r71 77 81 0.655813
r72 72 73 0.65228
r73 71 72 3.42052
r74 66 71 0.65409
r75 42 57 1.16709
r76 42 73 2.1395
r77 37 52 1.16709
r78 37 81 12.0712
r79 37 66 1.96931
r80 32 49 1.16709
r81 32 77 3.25093
r82 29 49 0.1
r83 21 57 0.50025
r84 18 52 0.50025
r85 8 21 4.37625
r86 6 18 4.37625
r87 4 29 0.123773
r88 2 29 0.123773
.ends

.subckt PM_G4_MAJ3_N3_AI 2 4 7 11 31 37 43 46 51 60 69 Vss
c43 69 Vss 4.20376e-19
c44 60 Vss 0.00685099f
c45 51 Vss 0.00640177f
c46 46 Vss 9.78141e-19
c47 43 Vss 0.00452529f
c48 37 Vss 0.12791f
c49 31 Vss 0.134433f
c50 7 Vss 1.43419f
c51 4 Vss 0.00143493f
r52 65 69 0.652036
r53 60 63 0.1
r54 51 63 1.16709
r55 51 69 13.7539
r56 46 65 3.501
r57 43 46 1.16709
r58 36 60 0.0238214
r59 36 37 2.334
r60 33 36 2.20433
r61 29 31 4.53833
r62 26 37 0.00605528
r63 25 31 0.00605528
r64 22 33 0.00605528
r65 21 29 0.00605528
r66 11 26 5.1348
r67 11 22 5.1348
r68 7 11 17.9718
r69 7 25 5.1348
r70 7 11 17.9718
r71 7 21 5.1348
r72 4 43 0.123773
r73 2 43 0.123773
.ends

.subckt PM_G4_MAJ3_N3_B 2 4 6 8 16 17 26 38 42 45 50 55 60 65 73 74 80 87 92 93
+ Vss
c63 93 Vss 4.8362e-19
c64 92 Vss 0.00212566f
c65 87 Vss 9.92513e-19
c66 80 Vss 6.85439e-19
c67 74 Vss 5.17886e-19
c68 73 Vss 0.00375307f
c69 65 Vss 0.00163151f
c70 60 Vss 0.00118605f
c71 55 Vss 0.00132948f
c72 50 Vss 0.00183658f
c73 45 Vss 7.01705e-19
c74 38 Vss 0.00124968f
c75 26 Vss 0.166484f
c76 20 Vss 0.0247918f
c77 17 Vss 0.0349747f
c78 16 Vss 0.185505f
c79 8 Vss 0.166484f
c80 4 Vss 0.180512f
c81 2 Vss 0.192541f
r82 91 93 0.65409
r83 91 92 3.42052
r84 87 92 0.65228
r85 83 87 2.1006
r86 80 83 2.04225
r87 73 80 0.0685365
r88 73 74 10.3363
r89 69 74 0.652036
r90 50 65 1.16709
r91 50 93 2.00578
r92 45 60 1.16709
r93 45 83 0.0416786
r94 38 55 1.16709
r95 38 69 1.66714
r96 38 42 0.0833571
r97 36 55 0.238214
r98 33 65 0.50025
r99 26 60 0.50025
r100 24 36 0.262036
r101 20 36 0.326018
r102 20 24 0.05835
r103 17 36 6.7686
r104 16 36 0.326018
r105 16 36 0.1167
r106 13 17 0.652036
r107 8 33 4.37625
r108 6 26 4.37625
r109 4 24 5.07645
r110 2 13 5.1348
.ends

.subckt PM_G4_MAJ3_N3_C 2 4 12 17 20 25 51 Vss
c18 25 Vss 0.0055264f
c19 20 Vss 6.62222e-19
c20 17 Vss 0.00968607f
c21 12 Vss 0.00811861f
r22 25 51 1.89637
r23 20 51 8.169
r24 17 25 1.16709
r25 12 20 1.16709
r26 4 17 0.123773
r27 2 12 0.123773
.ends

.subckt PM_G4_MAJ3_N3_Z 2 4 6 8 23 27 30 33 Vss
c31 30 Vss 0.00306612f
c32 27 Vss 0.00807893f
c33 23 Vss 0.00720868f
c34 8 Vss 0.00143493f
c35 6 Vss 0.00143493f
r36 33 35 11.4616
r37 30 33 1.37539
r38 27 35 1.16709
r39 23 30 1.16709
r40 8 27 0.123773
r41 6 23 0.123773
r42 4 27 0.123773
r43 2 23 0.123773
.ends

.subckt G4_MAJ3_N3  VDD VSS A B C Z
*
* Z	Z
* C	C
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI19.X0 N_BI_XI19.X0_D N_VSS_XI19.X0_PGD N_B_XI19.X0_CG N_VSS_XI19.X0_PGD
+ N_VDD_XI19.X0_S TIGFET_HPNW12
XI18.X0 N_AI_XI18.X0_D N_VSS_XI18.X0_PGD N_A_XI18.X0_CG N_VSS_XI18.X0_PGD
+ N_VDD_XI18.X0_S TIGFET_HPNW12
XI17.X0 N_BI_XI17.X0_D N_VDD_XI17.X0_PGD N_B_XI17.X0_CG N_VDD_XI17.X0_PGD
+ N_VSS_XI17.X0_S TIGFET_HPNW12
XI16.X0 N_AI_XI16.X0_D N_VDD_XI16.X0_PGD N_A_XI16.X0_CG N_VDD_XI16.X0_PGD
+ N_VSS_XI16.X0_S TIGFET_HPNW12
XI22.X0 N_Z_XI22.X0_D N_AI_XI22.X0_PGD N_BI_XI22.X0_CG N_AI_XI22.X0_PGD
+ N_A_XI22.X0_S TIGFET_HPNW12
XI21.X0 N_Z_XI21.X0_D N_AI_XI21.X0_PGD N_B_XI21.X0_CG N_AI_XI21.X0_PGD
+ N_C_XI21.X0_S TIGFET_HPNW12
XI23.X0 N_Z_XI23.X0_D N_A_XI23.X0_PGD N_B_XI23.X0_CG N_A_XI23.X0_PGD
+ N_A_XI23.X0_S TIGFET_HPNW12
XI20.X0 N_Z_XI20.X0_D N_A_XI20.X0_PGD N_BI_XI20.X0_CG N_A_XI20.X0_PGD
+ N_C_XI20.X0_S TIGFET_HPNW12
*
x_PM_G4_MAJ3_N3_VDD N_VDD_XI19.X0_S N_VDD_XI18.X0_S N_VDD_XI17.X0_PGD
+ N_VDD_XI16.X0_PGD N_VDD_c_62_p N_VDD_c_4_p N_VDD_c_74_p N_VDD_c_63_p
+ N_VDD_c_8_p N_VDD_c_55_p N_VDD_c_64_p N_VDD_c_6_p N_VDD_c_33_p N_VDD_c_3_p
+ N_VDD_c_5_p N_VDD_c_39_p N_VDD_c_38_p VDD N_VDD_c_40_p N_VDD_c_9_p
+ N_VDD_c_42_p N_VDD_c_13_p N_VDD_c_17_p N_VDD_c_35_p N_VDD_c_36_p N_VDD_c_14_p
+ N_VDD_c_18_p Vss PM_G4_MAJ3_N3_VDD
x_PM_G4_MAJ3_N3_VSS N_VSS_XI19.X0_PGD N_VSS_XI18.X0_PGD N_VSS_XI17.X0_S
+ N_VSS_XI16.X0_S N_VSS_c_80_n N_VSS_c_82_n N_VSS_c_84_n N_VSS_c_86_n
+ N_VSS_c_123_p N_VSS_c_125_p N_VSS_c_87_n N_VSS_c_91_n N_VSS_c_95_n
+ N_VSS_c_96_n N_VSS_c_99_n N_VSS_c_100_n N_VSS_c_104_n N_VSS_c_108_n
+ N_VSS_c_113_n N_VSS_c_115_n N_VSS_c_116_n N_VSS_c_118_n N_VSS_c_119_n
+ N_VSS_c_120_n N_VSS_c_121_n VSS Vss PM_G4_MAJ3_N3_VSS
x_PM_G4_MAJ3_N3_A N_A_XI18.X0_CG N_A_XI16.X0_CG N_A_XI22.X0_S N_A_XI23.X0_S
+ N_A_XI23.X0_PGD N_A_XI20.X0_PGD N_A_c_158_n N_A_c_193_p N_A_c_195_p
+ N_A_c_168_n N_A_c_219_p N_A_c_159_n A N_A_c_174_n N_A_c_163_n N_A_c_214_p
+ N_A_c_180_p N_A_c_222_p N_A_c_165_n N_A_c_206_p N_A_c_166_n N_A_c_207_p Vss
+ PM_G4_MAJ3_N3_A
x_PM_G4_MAJ3_N3_BI N_BI_XI19.X0_D N_BI_XI17.X0_D N_BI_XI22.X0_CG N_BI_XI20.X0_CG
+ N_BI_c_243_n N_BI_c_230_n N_BI_c_232_n N_BI_c_240_n N_BI_c_260_p N_BI_c_248_n
+ N_BI_c_249_n N_BI_c_250_n N_BI_c_271_p N_BI_c_274_p N_BI_c_251_n Vss
+ PM_G4_MAJ3_N3_BI
x_PM_G4_MAJ3_N3_AI N_AI_XI18.X0_D N_AI_XI16.X0_D N_AI_XI22.X0_PGD
+ N_AI_XI21.X0_PGD N_AI_c_290_n N_AI_c_291_n N_AI_c_292_n N_AI_c_295_n
+ N_AI_c_299_n N_AI_c_308_n N_AI_c_309_n Vss PM_G4_MAJ3_N3_AI
x_PM_G4_MAJ3_N3_B N_B_XI19.X0_CG N_B_XI17.X0_CG N_B_XI21.X0_CG N_B_XI23.X0_CG
+ N_B_c_332_n N_B_c_342_n N_B_c_380_n N_B_c_333_n B N_B_c_360_n N_B_c_345_n
+ N_B_c_348_n N_B_c_365_n N_B_c_350_n N_B_c_338_n N_B_c_356_n N_B_c_357_n
+ N_B_c_374_n N_B_c_377_n N_B_c_378_n Vss PM_G4_MAJ3_N3_B
x_PM_G4_MAJ3_N3_C N_C_XI21.X0_S N_C_XI20.X0_S N_C_c_394_n N_C_c_407_p
+ N_C_c_395_n N_C_c_397_n C Vss PM_G4_MAJ3_N3_C
x_PM_G4_MAJ3_N3_Z N_Z_XI22.X0_D N_Z_XI21.X0_D N_Z_XI23.X0_D N_Z_XI20.X0_D
+ N_Z_c_412_n N_Z_c_437_n N_Z_c_417_n Z Vss PM_G4_MAJ3_N3_Z
cc_1 N_VDD_XI17.X0_PGD N_VSS_XI19.X0_PGD 0.00200629f
cc_2 N_VDD_XI16.X0_PGD N_VSS_XI18.X0_PGD 0.00200315f
cc_3 N_VDD_c_3_p N_VSS_XI18.X0_PGD 3.80615e-19
cc_4 N_VDD_c_4_p N_VSS_c_80_n 0.00200629f
cc_5 N_VDD_c_5_p N_VSS_c_80_n 3.89167e-19
cc_6 N_VDD_c_6_p N_VSS_c_82_n 3.80615e-19
cc_7 N_VDD_c_5_p N_VSS_c_82_n 3.89167e-19
cc_8 N_VDD_c_8_p N_VSS_c_84_n 0.00200315f
cc_9 N_VDD_c_9_p N_VSS_c_84_n 3.00203e-19
cc_10 N_VDD_c_9_p N_VSS_c_86_n 3.89167e-19
cc_11 N_VDD_c_6_p N_VSS_c_87_n 4.35319e-19
cc_12 N_VDD_c_5_p N_VSS_c_87_n 0.00141228f
cc_13 N_VDD_c_13_p N_VSS_c_87_n 9.22325e-19
cc_14 N_VDD_c_14_p N_VSS_c_87_n 3.48267e-19
cc_15 N_VDD_c_3_p N_VSS_c_91_n 4.35319e-19
cc_16 N_VDD_c_9_p N_VSS_c_91_n 0.00141228f
cc_17 N_VDD_c_17_p N_VSS_c_91_n 8.59637e-19
cc_18 N_VDD_c_18_p N_VSS_c_91_n 3.48267e-19
cc_19 N_VDD_c_13_p N_VSS_c_95_n 8.49247e-19
cc_20 N_VDD_XI16.X0_PGD N_VSS_c_96_n 2.8629e-19
cc_21 N_VDD_c_17_p N_VSS_c_96_n 0.00515616f
cc_22 N_VDD_c_18_p N_VSS_c_96_n 9.58524e-19
cc_23 N_VDD_c_9_p N_VSS_c_99_n 0.00403878f
cc_24 N_VDD_c_6_p N_VSS_c_100_n 3.66936e-19
cc_25 N_VDD_c_5_p N_VSS_c_100_n 0.00114511f
cc_26 N_VDD_c_13_p N_VSS_c_100_n 3.99794e-19
cc_27 N_VDD_c_14_p N_VSS_c_100_n 6.489e-19
cc_28 N_VDD_c_3_p N_VSS_c_104_n 3.66936e-19
cc_29 N_VDD_c_9_p N_VSS_c_104_n 0.00114511f
cc_30 N_VDD_c_17_p N_VSS_c_104_n 3.99794e-19
cc_31 N_VDD_c_18_p N_VSS_c_104_n 6.489e-19
cc_32 N_VDD_c_6_p N_VSS_c_108_n 0.00412661f
cc_33 N_VDD_c_33_p N_VSS_c_108_n 0.00936637f
cc_34 N_VDD_c_3_p N_VSS_c_108_n 0.00380969f
cc_35 N_VDD_c_35_p N_VSS_c_108_n 0.00104624f
cc_36 N_VDD_c_36_p N_VSS_c_108_n 0.0010706f
cc_37 N_VDD_c_5_p N_VSS_c_113_n 0.00331675f
cc_38 N_VDD_c_38_p N_VSS_c_113_n 2.97469e-19
cc_39 N_VDD_c_39_p N_VSS_c_115_n 0.00106807f
cc_40 N_VDD_c_40_p N_VSS_c_116_n 2.97469e-19
cc_41 N_VDD_c_9_p N_VSS_c_116_n 0.00331675f
cc_42 N_VDD_c_42_p N_VSS_c_118_n 0.00106807f
cc_43 N_VDD_c_5_p N_VSS_c_119_n 0.00602033f
cc_44 N_VDD_c_5_p N_VSS_c_120_n 7.74609e-19
cc_45 N_VDD_c_9_p N_VSS_c_121_n 7.74609e-19
cc_46 N_VDD_XI16.X0_PGD N_A_c_158_n 3.96972e-19
cc_47 N_VDD_XI16.X0_PGD N_A_c_159_n 5.06189e-19
cc_48 N_VDD_c_9_p N_A_c_159_n 2.07512e-19
cc_49 N_VDD_c_17_p N_A_c_159_n 2.39252e-19
cc_50 N_VDD_c_18_p N_A_c_159_n 2.01254e-19
cc_51 N_VDD_c_13_p N_A_c_163_n 5.45323e-19
cc_52 N_VDD_c_14_p N_A_c_163_n 4.10732e-19
cc_53 N_VDD_c_33_p N_A_c_165_n 9.17955e-19
cc_54 N_VDD_c_33_p N_A_c_166_n 5.22471e-19
cc_55 N_VDD_c_55_p N_BI_c_230_n 3.43419e-19
cc_56 N_VDD_c_38_p N_BI_c_230_n 3.72199e-19
cc_57 N_VDD_c_55_p N_BI_c_232_n 3.48267e-19
cc_58 N_VDD_c_5_p N_BI_c_232_n 3.12875e-19
cc_59 N_VDD_c_38_p N_BI_c_232_n 5.2846e-19
cc_60 N_VDD_XI17.X0_PGD N_AI_XI22.X0_PGD 2.84861e-19
cc_61 N_VDD_XI16.X0_PGD N_AI_XI22.X0_PGD 3.10667e-19
cc_62 N_VDD_c_62_p N_AI_c_290_n 2.84861e-19
cc_63 N_VDD_c_63_p N_AI_c_291_n 3.10667e-19
cc_64 N_VDD_c_64_p N_AI_c_292_n 3.43419e-19
cc_65 N_VDD_c_40_p N_AI_c_292_n 3.72199e-19
cc_66 N_VDD_c_9_p N_AI_c_292_n 2.74986e-19
cc_67 N_VDD_c_64_p N_AI_c_295_n 3.48267e-19
cc_68 N_VDD_c_3_p N_AI_c_295_n 2.34601e-19
cc_69 N_VDD_c_40_p N_AI_c_295_n 5.226e-19
cc_70 N_VDD_c_9_p N_AI_c_295_n 2.9533e-19
cc_71 N_VDD_c_17_p N_AI_c_299_n 9.90259e-19
cc_72 N_VDD_c_33_p N_B_XI19.X0_CG 3.68219e-19
cc_73 N_VDD_XI17.X0_PGD N_B_c_332_n 4.01605e-19
cc_74 N_VDD_c_74_p N_B_c_333_n 2.01616e-19
cc_75 N_VDD_c_33_p N_B_c_333_n 3.58277e-19
cc_76 N_VDD_c_14_p N_B_c_333_n 2.07877e-19
cc_77 N_VSS_XI18.X0_PGD N_A_c_158_n 3.96972e-19
cc_78 N_VSS_c_123_p N_A_c_168_n 3.43419e-19
cc_79 N_VSS_c_123_p N_A_c_159_n 2.21087e-19
cc_80 N_VSS_c_125_p N_A_c_159_n 4.13509e-19
cc_81 N_VSS_c_95_n N_A_c_159_n 2.50981e-19
cc_82 N_VSS_c_96_n N_A_c_159_n 7.05313e-19
cc_83 N_VSS_c_99_n N_A_c_159_n 2.62883e-19
cc_84 N_VSS_c_123_p N_A_c_174_n 9.18655e-19
cc_85 N_VSS_c_95_n N_A_c_174_n 0.00202874f
cc_86 N_VSS_c_95_n N_A_c_163_n 0.00196507f
cc_87 N_VSS_c_104_n N_A_c_165_n 4.60155e-19
cc_88 N_VSS_c_108_n N_A_c_165_n 5.04162e-19
cc_89 N_VSS_c_91_n N_A_c_166_n 2.15082e-19
cc_90 N_VSS_c_123_p N_BI_c_230_n 3.43419e-19
cc_91 N_VSS_c_123_p N_BI_c_232_n 3.48267e-19
cc_92 N_VSS_c_95_n N_BI_c_232_n 0.00105024f
cc_93 N_VSS_c_108_n N_BI_c_232_n 0.00120568f
cc_94 N_VSS_c_119_n N_BI_c_232_n 2.38659e-19
cc_95 N_VSS_c_95_n N_BI_c_240_n 4.33962e-19
cc_96 N_VSS_c_119_n N_BI_c_240_n 6.35155e-19
cc_97 N_VSS_c_125_p N_AI_c_292_n 3.43419e-19
cc_98 N_VSS_c_96_n N_AI_c_292_n 3.48267e-19
cc_99 N_VSS_c_125_p N_AI_c_295_n 3.48267e-19
cc_100 N_VSS_c_91_n N_AI_c_295_n 0.00173332f
cc_101 N_VSS_c_96_n N_AI_c_295_n 0.00178201f
cc_102 N_VSS_c_108_n N_AI_c_295_n 0.00136931f
cc_103 N_VSS_c_96_n N_AI_c_299_n 0.00200998f
cc_104 N_VSS_c_99_n N_AI_c_299_n 0.00674978f
cc_105 N_VSS_c_96_n N_AI_c_308_n 2.82216e-19
cc_106 N_VSS_c_99_n N_AI_c_309_n 0.00178766f
cc_107 N_VSS_XI19.X0_PGD N_B_c_332_n 4.01605e-19
cc_108 N_VSS_c_108_n N_B_c_333_n 7.40204e-19
cc_109 N_VSS_c_95_n N_B_c_338_n 4.25717e-19
cc_110 N_VSS_c_125_p N_C_c_394_n 3.43419e-19
cc_111 N_VSS_c_125_p N_C_c_395_n 3.48267e-19
cc_112 N_VSS_c_96_n N_C_c_395_n 6.01757e-19
cc_113 N_A_c_180_p N_BI_XI22.X0_CG 2.10479e-19
cc_114 N_A_XI23.X0_PGD N_BI_c_243_n 9.65637e-19
cc_115 N_A_c_159_n N_BI_c_232_n 3.45962e-19
cc_116 N_A_c_174_n N_BI_c_232_n 5.71688e-19
cc_117 N_A_c_174_n N_BI_c_240_n 0.00169296f
cc_118 N_A_c_180_p N_BI_c_240_n 6.66847e-19
cc_119 N_A_c_174_n N_BI_c_248_n 3.37713e-19
cc_120 N_A_XI23.X0_PGD N_BI_c_249_n 0.00245019f
cc_121 N_A_c_180_p N_BI_c_250_n 9.24697e-19
cc_122 N_A_c_159_n N_BI_c_251_n 8.09947e-19
cc_123 N_A_XI23.X0_PGD N_AI_XI22.X0_PGD 0.0174035f
cc_124 N_A_c_174_n N_AI_XI22.X0_PGD 8.23587e-19
cc_125 N_A_c_180_p N_AI_XI22.X0_PGD 9.89767e-19
cc_126 N_A_c_193_p N_AI_c_290_n 0.00196311f
cc_127 N_A_c_180_p N_AI_c_290_n 0.00103585f
cc_128 N_A_c_195_p N_AI_c_291_n 0.00200674f
cc_129 N_A_c_158_n N_AI_c_292_n 6.90199e-19
cc_130 N_A_c_159_n N_AI_c_295_n 5.79974e-19
cc_131 N_A_c_159_n N_AI_c_299_n 0.00132412f
cc_132 N_A_XI23.X0_PGD N_B_XI23.X0_CG 9.65637e-19
cc_133 N_A_c_158_n N_B_c_332_n 0.0036037f
cc_134 N_A_c_159_n N_B_c_332_n 8.51862e-19
cc_135 N_A_c_166_n N_B_c_342_n 6.91203e-19
cc_136 N_A_c_159_n N_B_c_333_n 0.00120731f
cc_137 N_A_c_174_n N_B_c_333_n 0.00118668f
cc_138 N_A_c_180_p N_B_c_345_n 3.57869e-19
cc_139 N_A_c_206_p N_B_c_345_n 3.46877e-19
cc_140 N_A_c_207_p N_B_c_345_n 2.26741e-19
cc_141 N_A_c_159_n N_B_c_348_n 7.40468e-19
cc_142 N_A_c_174_n N_B_c_348_n 5.93411e-19
cc_143 N_A_XI23.X0_PGD N_B_c_350_n 0.00312702f
cc_144 N_A_c_206_p N_B_c_350_n 2.30774e-19
cc_145 N_A_c_159_n N_B_c_338_n 0.00230073f
cc_146 N_A_c_174_n N_B_c_338_n 0.00203212f
cc_147 N_A_c_214_p N_B_c_338_n 3.55185e-19
cc_148 N_A_c_180_p N_B_c_338_n 4.84888e-19
cc_149 N_A_c_159_n N_B_c_356_n 4.20277e-19
cc_150 N_A_c_159_n N_B_c_357_n 2.29222e-19
cc_151 N_A_c_168_n N_Z_c_412_n 3.43419e-19
cc_152 N_A_c_219_p N_Z_c_412_n 3.43419e-19
cc_153 N_A_c_214_p N_Z_c_412_n 3.48267e-19
cc_154 N_A_c_180_p N_Z_c_412_n 5.52794e-19
cc_155 N_A_c_222_p N_Z_c_412_n 3.48267e-19
cc_156 N_A_XI23.X0_PGD N_Z_c_417_n 6.68421e-19
cc_157 N_A_c_168_n N_Z_c_417_n 3.48267e-19
cc_158 N_A_c_219_p N_Z_c_417_n 3.48267e-19
cc_159 N_A_c_174_n N_Z_c_417_n 0.00158522f
cc_160 N_A_c_214_p N_Z_c_417_n 7.9714e-19
cc_161 N_A_c_180_p N_Z_c_417_n 9.31302e-19
cc_162 N_A_c_222_p N_Z_c_417_n 8.16241e-19
cc_163 N_BI_XI22.X0_CG N_AI_XI22.X0_PGD 9.47088e-19
cc_164 N_BI_c_248_n N_AI_XI22.X0_PGD 0.00312702f
cc_165 N_BI_c_251_n N_AI_c_295_n 2.92168e-19
cc_166 N_BI_c_240_n N_AI_c_299_n 3.11073e-19
cc_167 N_BI_c_230_n N_B_c_332_n 6.90199e-19
cc_168 N_BI_c_240_n N_B_c_333_n 0.0014575f
cc_169 N_BI_c_240_n N_B_c_360_n 6.83975e-19
cc_170 N_BI_c_248_n N_B_c_360_n 4.99367e-19
cc_171 N_BI_c_260_p N_B_c_345_n 0.0018485f
cc_172 N_BI_c_249_n N_B_c_345_n 4.99367e-19
cc_173 N_BI_c_250_n N_B_c_345_n 0.00165504f
cc_174 N_BI_c_248_n N_B_c_365_n 0.00521054f
cc_175 N_BI_c_249_n N_B_c_365_n 7.2092e-19
cc_176 N_BI_c_260_p N_B_c_350_n 4.99367e-19
cc_177 N_BI_c_248_n N_B_c_350_n 6.22265e-19
cc_178 N_BI_c_249_n N_B_c_350_n 0.00494884f
cc_179 N_BI_c_240_n N_B_c_338_n 0.00536154f
cc_180 N_BI_c_240_n N_B_c_357_n 2.67017e-19
cc_181 N_BI_c_250_n N_B_c_357_n 0.0013533f
cc_182 N_BI_c_271_p N_B_c_357_n 0.00340518f
cc_183 N_BI_c_240_n N_B_c_374_n 4.99817e-19
cc_184 N_BI_c_250_n N_B_c_374_n 9.84686e-19
cc_185 N_BI_c_274_p N_B_c_374_n 7.60478e-19
cc_186 N_BI_c_271_p N_B_c_377_n 0.00181541f
cc_187 N_BI_c_240_n N_B_c_378_n 0.00145553f
cc_188 N_BI_c_250_n N_B_c_378_n 8.77567e-19
cc_189 N_BI_c_240_n N_C_c_397_n 9.46412e-19
cc_190 N_BI_c_260_p N_C_c_397_n 0.00112215f
cc_191 N_BI_c_274_p N_C_c_397_n 2.41224e-19
cc_192 N_BI_c_240_n N_Z_c_417_n 0.00190811f
cc_193 N_BI_c_260_p N_Z_c_417_n 0.00192905f
cc_194 N_BI_c_248_n N_Z_c_417_n 8.66889e-19
cc_195 N_BI_c_249_n N_Z_c_417_n 8.66889e-19
cc_196 N_BI_c_250_n N_Z_c_417_n 0.00108781f
cc_197 N_BI_c_271_p N_Z_c_417_n 0.00210701f
cc_198 N_BI_c_274_p N_Z_c_417_n 0.00102097f
cc_199 N_AI_XI22.X0_PGD N_B_c_380_n 9.65637e-19
cc_200 N_AI_c_299_n N_B_c_360_n 3.12862e-19
cc_201 N_AI_c_308_n N_B_c_360_n 2.26741e-19
cc_202 N_AI_XI22.X0_PGD N_B_c_365_n 0.00312702f
cc_203 N_AI_c_299_n N_B_c_338_n 0.00252591f
cc_204 N_AI_c_299_n N_C_c_395_n 0.00111024f
cc_205 N_AI_c_299_n N_C_c_397_n 0.0016345f
cc_206 N_AI_XI22.X0_PGD N_Z_c_417_n 3.73496e-19
cc_207 N_B_c_338_n N_C_c_395_n 4.14759e-19
cc_208 N_B_c_345_n N_C_c_397_n 8.23684e-19
cc_209 N_B_c_338_n N_C_c_397_n 3.71981e-19
cc_210 N_B_c_374_n N_C_c_397_n 0.0032187f
cc_211 N_B_c_360_n N_Z_c_417_n 0.00192136f
cc_212 N_B_c_345_n N_Z_c_417_n 0.0019232f
cc_213 N_B_c_365_n N_Z_c_417_n 8.66889e-19
cc_214 N_B_c_350_n N_Z_c_417_n 8.66889e-19
cc_215 N_B_c_357_n N_Z_c_417_n 4.75654e-19
cc_216 N_C_c_394_n N_Z_c_437_n 3.43419e-19
cc_217 N_C_c_407_p N_Z_c_437_n 3.43419e-19
cc_218 N_C_c_395_n N_Z_c_437_n 3.48267e-19
cc_219 N_C_c_397_n N_Z_c_437_n 3.48267e-19
cc_220 N_C_c_395_n N_Z_c_417_n 6.20216e-19
cc_221 N_C_c_397_n N_Z_c_417_n 0.00134739f
*
.ends
*
*
.subckt MAJ3_HPNW12 A B C Y VDD VSS
xgate (VDD VSS A B C Y) G4_MAJ3_N3
.ends
*
* File: G3_MIN3_T6_N3.pex.netlist
* Created: Mon Apr  4 15:49:45 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MIN3_T6_N3_VSS 2 4 6 8 10 12 27 32 37 40 42 45 53 57 60 65 70 75
+ 88 89 93 99 101 106 109 Vss
c64 107 Vss 6.47574e-19
c65 106 Vss 0.00464148f
c66 101 Vss 0.00213175f
c67 99 Vss 0.0082833f
c68 94 Vss 0.00138375f
c69 93 Vss 0.00819383f
c70 89 Vss 6.61473e-19
c71 88 Vss 0.0060976f
c72 75 Vss 0.006288f
c73 70 Vss 1.73335e-19
c74 65 Vss 0.00209248f
c75 60 Vss 0.00138481f
c76 57 Vss 0.0103194f
c77 53 Vss 0.00454903f
c78 45 Vss 0.0856842f
c79 42 Vss 0.0855647f
c80 37 Vss 0.0648277f
c81 32 Vss 0.103906f
c82 27 Vss 0.306999f
c83 22 Vss 0.141041f
c84 10 Vss 0.186558f
c85 8 Vss 0.00171982f
c86 6 Vss 0.188337f
c87 2 Vss 0.185627f
r88 106 109 0.326018
r89 105 106 5.50157
r90 101 105 0.655813
r91 100 107 0.494161
r92 99 109 0.326018
r93 99 100 13.0037
r94 95 107 0.128424
r95 93 107 0.494161
r96 93 94 10.0862
r97 88 94 0.652036
r98 87 89 0.655813
r99 87 88 16.4214
r100 70 101 1.82344
r101 65 95 6.16843
r102 60 75 1.16709
r103 60 89 1.82344
r104 57 70 1.16709
r105 53 65 1.16709
r106 45 47 1.8672
r107 42 44 1.8672
r108 40 75 0.50025
r109 37 40 1.92555
r110 33 47 0.0685365
r111 32 34 0.652036
r112 32 33 2.8008
r113 29 47 0.5835
r114 28 42 0.0685365
r115 27 45 0.0685365
r116 27 28 10.9698
r117 24 44 0.5835
r118 23 37 0.0685365
r119 22 44 0.0685365
r120 22 23 4.7847
r121 12 57 0.123773
r122 10 34 5.1348
r123 8 53 0.123773
r124 6 29 5.1348
r125 4 53 0.123773
r126 2 24 5.1348
.ends

.subckt PM_G3_MIN3_T6_N3_VDD 2 4 6 8 10 12 27 32 42 45 53 57 60 61 63 65 69 71
+ 73 78 81 83 Vss
c74 83 Vss 0.00747336f
c75 79 Vss 7.84502e-19
c76 78 Vss 0.00603664f
c77 73 Vss 0.00149586f
c78 71 Vss 0.0125181f
c79 69 Vss 0.00223179f
c80 65 Vss 0.00180228f
c81 63 Vss 7.51405e-19
c82 62 Vss 0.00180268f
c83 61 Vss 0.00800879f
c84 60 Vss 0.00954496f
c85 57 Vss 0.00979559f
c86 53 Vss 0.00450493f
c87 45 Vss 0.0849231f
c88 42 Vss 0.0854945f
c89 38 Vss 0.0711342f
c90 32 Vss 0.106731f
c91 27 Vss 0.308123f
c92 22 Vss 0.144485f
c93 12 Vss 0.187032f
c94 8 Vss 0.187847f
c95 6 Vss 0.00171982f
c96 4 Vss 0.18764f
r97 78 81 0.349767
r98 77 78 5.50157
r99 73 81 0.306046
r100 73 75 1.82344
r101 72 79 0.494161
r102 71 77 0.652036
r103 71 72 13.0037
r104 67 79 0.128424
r105 67 69 6.16843
r106 65 83 1.16709
r107 63 65 1.82344
r108 61 79 0.494161
r109 61 62 10.0862
r110 60 63 0.655813
r111 59 62 0.652036
r112 59 60 16.4214
r113 57 75 1.16709
r114 53 69 1.16709
r115 45 46 1.8672
r116 42 43 1.8672
r117 38 83 0.50025
r118 38 40 1.92555
r119 33 45 0.0685365
r120 32 34 0.652036
r121 32 33 2.8008
r122 29 45 0.5835
r123 28 43 0.0685365
r124 27 46 0.0685365
r125 27 28 10.9698
r126 24 42 0.5835
r127 23 40 0.0685365
r128 22 42 0.0685365
r129 22 23 4.7847
r130 12 34 5.1348
r131 10 57 0.123773
r132 8 29 5.1348
r133 6 53 0.123773
r134 4 24 5.1348
r135 2 53 0.123773
.ends

.subckt PM_G3_MIN3_T6_N3_Z 2 4 6 8 10 12 32 36 41 45 49 53 55 59 63 67 Vss
c55 67 Vss 3.51451e-19
c56 65 Vss 2.45386e-19
c57 63 Vss 0.00102688f
c58 59 Vss 7.58182e-19
c59 55 Vss 0.0050105f
c60 53 Vss 6.51205e-19
c61 49 Vss 5.16244e-19
c62 45 Vss 0.00816234f
c63 41 Vss 0.00751221f
c64 36 Vss 0.00857712f
c65 32 Vss 0.00789336f
c66 12 Vss 0.00171982f
c67 10 Vss 0.00171982f
r68 61 67 0.494161
r69 61 63 3.95946
r70 57 67 0.494161
r71 57 59 3.95946
r72 56 65 0.128424
r73 55 67 0.128424
r74 55 56 10.3363
r75 51 65 0.494161
r76 51 53 3.95946
r77 47 65 0.494161
r78 47 49 3.95946
r79 45 63 1.16709
r80 41 59 1.16709
r81 36 53 1.16709
r82 32 49 1.16709
r83 12 45 0.123773
r84 10 41 0.123773
r85 8 45 0.123773
r86 6 41 0.123773
r87 4 36 0.123773
r88 2 32 0.123773
.ends

.subckt PM_G3_MIN3_T6_N3_C 2 4 6 8 14 20 26 33 38 43 Vss
c33 43 Vss 0.00462472f
c34 38 Vss 0.00103857f
c35 33 Vss 0.00642701f
c36 26 Vss 7.12876e-22
c37 20 Vss 0.486644f
c38 14 Vss 0.489687f
r39 33 43 1.16709
r40 29 38 1.16709
r41 29 33 11.5033
r42 26 29 0.166714
r43 20 43 0.50025
r44 14 38 0.50025
r45 6 8 12.7203
r46 6 20 4.37625
r47 2 4 12.7203
r48 2 14 4.37625
.ends

.subckt PM_G3_MIN3_T6_N3_B 2 4 6 8 17 18 26 29 32 35 Vss
c31 35 Vss 0.00167659f
c32 26 Vss 0.0837857f
c33 18 Vss 0.034641f
c34 17 Vss 0.09638f
c35 6 Vss 0.506992f
c36 2 Vss 0.554218f
r37 32 35 1.16709
r38 29 32 0.0729375
r39 24 35 0.0476429
r40 24 26 1.92555
r41 17 19 0.652036
r42 17 18 2.8008
r43 14 26 0.0685365
r44 13 18 0.652036
r45 6 8 12.7203
r46 6 19 5.1348
r47 4 14 5.1348
r48 2 4 12.7203
r49 2 13 5.1348
.ends

.subckt PM_G3_MIN3_T6_N3_A 2 4 6 8 17 29 34 38 41 46 Vss
c29 46 Vss 0.00528506f
c30 41 Vss 0.00159958f
c31 38 Vss 3.66482e-19
c32 34 Vss 0.00172621f
c33 29 Vss 3.54075e-22
c34 26 Vss 0.0871371f
c35 6 Vss 0.515115f
c36 2 Vss 0.485149f
r37 34 46 1.16709
r38 34 38 0.109406
r39 29 41 1.16709
r40 29 34 5.03269
r41 24 46 0.0476429
r42 24 26 1.92555
r43 19 26 0.0685365
r44 17 41 0.50025
r45 8 19 5.1348
r46 6 8 12.7203
r47 4 17 4.37625
r48 2 4 12.7203
.ends

.subckt G3_MIN3_T6_N3  VSS VDD Z C B A
*
* A	A
* B	B
* C	C
* Z	Z
* VDD	VDD
* VSS	VSS
XI24.X0 N_Z_XI24.X0_D N_VSS_XI24.X0_PGD N_C_XI24.X0_CG N_B_XI24.X0_PGS
+ N_VDD_XI24.X0_S TIGFET_HPNW12
XI20.X0 N_Z_XI20.X0_D N_VDD_XI20.X0_PGD N_C_XI20.X0_CG N_B_XI20.X0_PGS
+ N_VSS_XI20.X0_S TIGFET_HPNW12
XI23.X0 N_Z_XI23.X0_D N_VSS_XI23.X0_PGD N_A_XI23.X0_CG N_B_XI23.X0_PGS
+ N_VDD_XI23.X0_S TIGFET_HPNW12
XI22.X0 N_Z_XI22.X0_D N_VDD_XI22.X0_PGD N_A_XI22.X0_CG N_B_XI22.X0_PGS
+ N_VSS_XI22.X0_S TIGFET_HPNW12
XI25.X0 N_Z_XI25.X0_D N_VSS_XI25.X0_PGD N_C_XI25.X0_CG N_A_XI25.X0_PGS
+ N_VDD_XI25.X0_S TIGFET_HPNW12
XI21.X0 N_Z_XI21.X0_D N_VDD_XI21.X0_PGD N_C_XI21.X0_CG N_A_XI21.X0_PGS
+ N_VSS_XI21.X0_S TIGFET_HPNW12
*
x_PM_G3_MIN3_T6_N3_VSS N_VSS_XI24.X0_PGD N_VSS_XI20.X0_S N_VSS_XI23.X0_PGD
+ N_VSS_XI22.X0_S N_VSS_XI25.X0_PGD N_VSS_XI21.X0_S N_VSS_c_19_p N_VSS_c_22_p
+ N_VSS_c_6_p N_VSS_c_12_p N_VSS_c_13_p N_VSS_c_46_p N_VSS_c_4_p N_VSS_c_29_p
+ N_VSS_c_7_p N_VSS_c_17_p N_VSS_c_23_p N_VSS_c_8_p N_VSS_c_9_p N_VSS_c_10_p
+ N_VSS_c_18_p N_VSS_c_43_p N_VSS_c_24_p N_VSS_c_62_p VSS Vss
+ PM_G3_MIN3_T6_N3_VSS
x_PM_G3_MIN3_T6_N3_VDD N_VDD_XI24.X0_S N_VDD_XI20.X0_PGD N_VDD_XI23.X0_S
+ N_VDD_XI22.X0_PGD N_VDD_XI25.X0_S N_VDD_XI21.X0_PGD N_VDD_c_68_n N_VDD_c_137_p
+ N_VDD_c_130_p N_VDD_c_129_p N_VDD_c_69_n N_VDD_c_96_p N_VDD_c_70_n
+ N_VDD_c_75_n N_VDD_c_79_n N_VDD_c_80_n N_VDD_c_83_n N_VDD_c_85_n N_VDD_c_87_n
+ N_VDD_c_119_p VDD N_VDD_c_89_n Vss PM_G3_MIN3_T6_N3_VDD
x_PM_G3_MIN3_T6_N3_Z N_Z_XI24.X0_D N_Z_XI20.X0_D N_Z_XI23.X0_D N_Z_XI22.X0_D
+ N_Z_XI25.X0_D N_Z_XI21.X0_D N_Z_c_154_n N_Z_c_139_n N_Z_c_159_n N_Z_c_141_n
+ N_Z_c_145_n N_Z_c_146_n N_Z_c_149_n N_Z_c_172_n N_Z_c_151_n Z Vss
+ PM_G3_MIN3_T6_N3_Z
x_PM_G3_MIN3_T6_N3_C N_C_XI24.X0_CG N_C_XI20.X0_CG N_C_XI25.X0_CG N_C_XI21.X0_CG
+ N_C_c_194_n N_C_c_195_n C N_C_c_196_n N_C_c_197_n N_C_c_198_n Vss
+ PM_G3_MIN3_T6_N3_C
x_PM_G3_MIN3_T6_N3_B N_B_XI24.X0_PGS N_B_XI20.X0_PGS N_B_XI23.X0_PGS
+ N_B_XI22.X0_PGS N_B_c_231_n N_B_c_232_n N_B_c_240_n B N_B_c_234_n N_B_c_242_n
+ Vss PM_G3_MIN3_T6_N3_B
x_PM_G3_MIN3_T6_N3_A N_A_XI23.X0_CG N_A_XI22.X0_CG N_A_XI25.X0_PGS
+ N_A_XI21.X0_PGS N_A_c_274_n N_A_c_259_n N_A_c_261_n A N_A_c_269_n N_A_c_270_n
+ Vss PM_G3_MIN3_T6_N3_A
cc_1 N_VSS_XI24.X0_PGD N_VDD_XI20.X0_PGD 6.54383e-19
cc_2 N_VSS_XI23.X0_PGD N_VDD_XI22.X0_PGD 6.54383e-19
cc_3 N_VSS_XI25.X0_PGD N_VDD_XI21.X0_PGD 6.43556e-19
cc_4 N_VSS_c_4_p N_VDD_c_68_n 5.08814e-19
cc_5 N_VSS_c_4_p N_VDD_c_69_n 7.73686e-19
cc_6 N_VSS_c_6_p N_VDD_c_70_n 2.63314e-19
cc_7 N_VSS_c_7_p N_VDD_c_70_n 0.00161042f
cc_8 N_VSS_c_8_p N_VDD_c_70_n 0.00115993f
cc_9 N_VSS_c_9_p N_VDD_c_70_n 0.00777883f
cc_10 N_VSS_c_10_p N_VDD_c_70_n 0.00186982f
cc_11 N_VSS_c_6_p N_VDD_c_75_n 8.77582e-19
cc_12 N_VSS_c_12_p N_VDD_c_75_n 3.72495e-19
cc_13 N_VSS_c_13_p N_VDD_c_75_n 7.64639e-19
cc_14 N_VSS_c_7_p N_VDD_c_75_n 9.97468e-19
cc_15 N_VSS_c_9_p N_VDD_c_79_n 0.00179061f
cc_16 N_VSS_c_7_p N_VDD_c_80_n 3.76254e-19
cc_17 N_VSS_c_17_p N_VDD_c_80_n 2.77394e-19
cc_18 N_VSS_c_18_p N_VDD_c_80_n 4.66156e-19
cc_19 N_VSS_c_19_p N_VDD_c_83_n 0.00120485f
cc_20 N_VSS_c_7_p N_VDD_c_83_n 4.38149e-19
cc_21 N_VSS_c_19_p N_VDD_c_85_n 8.70027e-19
cc_22 N_VSS_c_22_p N_VDD_c_85_n 8.24361e-19
cc_23 N_VSS_c_23_p N_VDD_c_87_n 2.543e-19
cc_24 N_VSS_c_24_p N_VDD_c_87_n 0.00120656f
cc_25 N_VSS_c_8_p N_VDD_c_89_n 2.36483e-19
cc_26 N_VSS_c_4_p N_Z_c_139_n 3.43419e-19
cc_27 N_VSS_c_17_p N_Z_c_139_n 3.48267e-19
cc_28 N_VSS_c_4_p N_Z_c_141_n 3.43419e-19
cc_29 N_VSS_c_29_p N_Z_c_141_n 3.43419e-19
cc_30 N_VSS_c_17_p N_Z_c_141_n 3.48267e-19
cc_31 N_VSS_c_23_p N_Z_c_141_n 3.48267e-19
cc_32 N_VSS_c_9_p N_Z_c_145_n 0.00213783f
cc_33 N_VSS_c_4_p N_Z_c_146_n 3.48267e-19
cc_34 N_VSS_c_17_p N_Z_c_146_n 5.02484e-19
cc_35 N_VSS_c_18_p N_Z_c_146_n 4.85461e-19
cc_36 N_VSS_c_4_p N_Z_c_149_n 4.81023e-19
cc_37 N_VSS_c_17_p N_Z_c_149_n 6.34336e-19
cc_38 N_VSS_c_29_p N_Z_c_151_n 3.48267e-19
cc_39 N_VSS_c_17_p N_Z_c_151_n 5.37696e-19
cc_40 N_VSS_c_23_p N_Z_c_151_n 5.71987e-19
cc_41 N_VSS_XI24.X0_PGD N_C_c_194_n 4.30517e-19
cc_42 N_VSS_XI25.X0_PGD N_C_c_195_n 4.94554e-19
cc_43 N_VSS_c_43_p N_C_c_196_n 5.18193e-19
cc_44 N_VSS_XI24.X0_PGD N_C_c_197_n 4.3583e-19
cc_45 N_VSS_XI25.X0_PGD N_C_c_198_n 3.76133e-19
cc_46 N_VSS_c_46_p N_C_c_198_n 2.17009e-19
cc_47 N_VSS_XI24.X0_PGD N_B_XI24.X0_PGS 0.00109504f
cc_48 N_VSS_XI23.X0_PGD N_B_XI24.X0_PGS 2.15671e-19
cc_49 N_VSS_XI23.X0_PGD N_B_XI23.X0_PGS 0.00177732f
cc_50 N_VSS_XI25.X0_PGD N_B_XI23.X0_PGS 2.22194e-19
cc_51 N_VSS_c_46_p N_B_c_231_n 0.00177732f
cc_52 N_VSS_c_19_p N_B_c_232_n 0.00722404f
cc_53 N_VSS_c_13_p N_B_c_232_n 0.00109504f
cc_54 N_VSS_c_17_p N_B_c_234_n 2.11465e-19
cc_55 N_VSS_c_9_p N_B_c_234_n 2.74582e-19
cc_56 N_VSS_c_18_p N_B_c_234_n 4.28832e-19
cc_57 N_VSS_c_19_p N_A_XI23.X0_CG 2.64949e-19
cc_58 N_VSS_c_17_p N_A_c_259_n 3.13396e-19
cc_59 N_VSS_c_43_p N_A_c_259_n 5.88825e-19
cc_60 N_VSS_c_17_p N_A_c_261_n 0.00159318f
cc_61 N_VSS_c_43_p N_A_c_261_n 0.00925582f
cc_62 N_VSS_c_62_p N_A_c_261_n 7.74234e-19
cc_63 N_VSS_c_43_p A 5.88825e-19
cc_64 N_VSS_c_62_p A 3.28646e-19
cc_65 N_VDD_c_69_n N_Z_c_154_n 3.43419e-19
cc_66 N_VDD_c_70_n N_Z_c_154_n 3.70842e-19
cc_67 N_VDD_c_75_n N_Z_c_154_n 2.74986e-19
cc_68 N_VDD_c_83_n N_Z_c_154_n 3.48267e-19
cc_69 N_VDD_c_70_n N_Z_c_139_n 3.70842e-19
cc_70 N_VDD_c_69_n N_Z_c_159_n 3.43419e-19
cc_71 N_VDD_c_96_p N_Z_c_159_n 3.43419e-19
cc_72 N_VDD_c_83_n N_Z_c_159_n 3.48267e-19
cc_73 N_VDD_c_85_n N_Z_c_159_n 2.74986e-19
cc_74 N_VDD_c_87_n N_Z_c_159_n 3.72199e-19
cc_75 N_VDD_c_69_n N_Z_c_145_n 3.48267e-19
cc_76 N_VDD_c_70_n N_Z_c_145_n 0.00440367f
cc_77 N_VDD_c_75_n N_Z_c_145_n 5.29921e-19
cc_78 N_VDD_c_83_n N_Z_c_145_n 7.15874e-19
cc_79 N_VDD_c_69_n N_Z_c_149_n 4.81023e-19
cc_80 N_VDD_c_75_n N_Z_c_149_n 3.00455e-19
cc_81 N_VDD_c_83_n N_Z_c_149_n 8.48441e-19
cc_82 N_VDD_c_85_n N_Z_c_149_n 4.56827e-19
cc_83 N_VDD_c_69_n N_Z_c_172_n 3.48267e-19
cc_84 N_VDD_c_96_p N_Z_c_172_n 3.48267e-19
cc_85 N_VDD_c_83_n N_Z_c_172_n 7.23486e-19
cc_86 N_VDD_c_85_n N_Z_c_172_n 4.06373e-19
cc_87 N_VDD_c_87_n N_Z_c_172_n 8.5731e-19
cc_88 N_VDD_c_70_n C 2.30446e-19
cc_89 N_VDD_c_75_n C 0.00138543f
cc_90 N_VDD_c_83_n C 0.00115642f
cc_91 N_VDD_c_75_n N_C_c_196_n 7.64872e-19
cc_92 N_VDD_c_83_n N_C_c_196_n 0.00221688f
cc_93 N_VDD_c_85_n N_C_c_196_n 0.0053512f
cc_94 N_VDD_c_119_p N_C_c_196_n 6.92542e-19
cc_95 N_VDD_c_75_n N_C_c_197_n 4.58746e-19
cc_96 N_VDD_c_83_n N_C_c_197_n 8.66889e-19
cc_97 N_VDD_c_83_n N_C_c_198_n 2.22969e-19
cc_98 N_VDD_c_85_n N_C_c_198_n 2.64043e-19
cc_99 N_VDD_c_119_p N_C_c_198_n 4.74797e-19
cc_100 N_VDD_XI20.X0_PGD N_B_XI24.X0_PGS 0.00135245f
cc_101 N_VDD_XI22.X0_PGD N_B_XI24.X0_PGS 4.12959e-19
cc_102 N_VDD_c_68_n N_B_XI23.X0_PGS 0.00108553f
cc_103 N_VDD_c_68_n N_B_c_240_n 0.00256877f
cc_104 N_VDD_c_129_p N_B_c_240_n 4.12959e-19
cc_105 N_VDD_c_130_p N_B_c_242_n 0.00495207f
cc_106 N_VDD_c_89_n N_B_c_242_n 4.60491e-19
cc_107 N_VDD_XI22.X0_PGD N_A_XI23.X0_CG 4.83278e-19
cc_108 N_VDD_XI21.X0_PGD N_A_XI25.X0_PGS 0.00150004f
cc_109 N_VDD_c_85_n N_A_XI25.X0_PGS 2.05774e-19
cc_110 N_VDD_XI22.X0_PGD N_A_c_269_n 5.50272e-19
cc_111 N_VDD_XI21.X0_PGD N_A_c_270_n 3.23173e-19
cc_112 N_VDD_c_137_p N_A_c_270_n 0.00145458f
cc_113 N_VDD_c_129_p N_A_c_270_n 2.17009e-19
cc_114 N_Z_c_145_n N_C_c_194_n 2.87038e-19
cc_115 N_Z_c_146_n N_C_c_194_n 2.87038e-19
cc_116 N_Z_c_149_n N_C_c_194_n 7.3418e-19
cc_117 N_Z_c_172_n N_C_c_195_n 0.00103972f
cc_118 N_Z_c_149_n C 2.05514e-19
cc_119 N_Z_c_149_n N_C_c_196_n 0.00135375f
cc_120 N_Z_c_172_n N_C_c_196_n 2.38669e-19
cc_121 N_Z_c_149_n N_C_c_197_n 2.28309e-19
cc_122 N_Z_c_149_n N_B_XI24.X0_PGS 7.69255e-19
cc_123 N_Z_c_149_n N_B_XI23.X0_PGS 8.11898e-19
cc_124 N_Z_c_149_n N_B_c_234_n 2.98201e-19
cc_125 N_Z_c_149_n N_B_c_242_n 2.18216e-19
cc_126 N_Z_c_149_n N_A_XI23.X0_CG 7.49661e-19
cc_127 N_Z_c_149_n N_A_c_274_n 2.18216e-19
cc_128 N_Z_c_149_n N_A_c_259_n 2.14102e-19
cc_129 N_Z_c_149_n N_A_c_261_n 2.49841e-19
cc_130 N_Z_c_151_n N_A_c_261_n 4.09814e-19
cc_131 N_C_c_194_n N_B_XI24.X0_PGS 0.00849032f
cc_132 N_C_c_197_n N_B_XI24.X0_PGS 3.76133e-19
cc_133 N_C_c_194_n N_B_XI23.X0_PGS 6.67601e-19
cc_134 N_C_c_195_n N_B_XI23.X0_PGS 4.29907e-19
cc_135 N_C_c_195_n N_A_XI23.X0_CG 0.00200107f
cc_136 N_C_c_195_n N_A_XI25.X0_PGS 0.00801113f
cc_137 N_C_c_196_n N_A_c_261_n 0.00114292f
cc_138 N_B_XI24.X0_PGS N_A_XI23.X0_CG 8.40291e-19
cc_139 N_B_XI23.X0_PGS N_A_XI23.X0_CG 0.00774979f
cc_140 N_B_c_234_n N_A_c_259_n 3.39698e-19
cc_141 N_B_c_242_n N_A_c_259_n 3.48267e-19
cc_142 N_B_c_234_n N_A_c_269_n 3.48267e-19
cc_143 N_B_c_242_n N_A_c_269_n 5.15124e-19
*
.ends
*
*
.subckt MIN3_HPNW12 A B C Y VDD VSS
xgate (VSS VDD Y C B A) G3_MIN3_T6_N3
.ends
*
* File: G4_MUX2_N3.pex.netlist
* Created: Tue Mar 15 11:34:09 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MUX2_N3_VDD 2 4 6 8 10 12 14 16 18 20 38 49 51 58 64 72 77 81 84
+ 85 89 93 95 96 99 101 105 107 111 113 115 120 122 124 125 126 127 128 134 139
+ 148 Vss
c131 148 Vss 0.00702165f
c132 139 Vss 0.00462928f
c133 134 Vss 0.00483792f
c134 128 Vss 4.52364e-19
c135 127 Vss 2.39889e-19
c136 126 Vss 4.24532e-19
c137 125 Vss 2.39889e-19
c138 122 Vss 0.00282332f
c139 120 Vss 0.0106931f
c140 115 Vss 0.00186946f
c141 113 Vss 0.006422f
c142 111 Vss 8.80889e-19
c143 107 Vss 0.00804399f
c144 105 Vss 0.00134677f
c145 101 Vss 0.00193004f
c146 99 Vss 3.98903e-19
c147 96 Vss 6.1175e-19
c148 95 Vss 0.00358057f
c149 93 Vss 0.00108621f
c150 89 Vss 0.00158874f
c151 86 Vss 0.00176185f
c152 85 Vss 0.0067647f
c153 84 Vss 0.00573691f
c154 81 Vss 0.00850511f
c155 77 Vss 0.00688835f
c156 72 Vss 0.00820121f
c157 64 Vss 8.40042e-20
c158 59 Vss 0.0806024f
c159 58 Vss 0.103898f
c160 49 Vss 0.0356247f
c161 48 Vss 0.101315f
c162 39 Vss 0.0367394f
c163 38 Vss 0.101469f
c164 18 Vss 0.188795f
c165 16 Vss 0.00143493f
c166 14 Vss 0.191141f
c167 10 Vss 0.187414f
c168 8 Vss 0.189706f
c169 6 Vss 0.190935f
c170 4 Vss 0.189249f
r171 121 128 0.551426
r172 121 122 5.50157
r173 120 128 0.551426
r174 119 120 18.3386
r175 115 128 0.0828784
r176 115 117 1.82344
r177 114 127 0.494161
r178 113 119 0.652036
r179 113 114 10.1279
r180 111 148 1.16709
r181 109 127 0.128424
r182 109 111 2.16729
r183 108 126 0.494161
r184 107 122 0.652036
r185 107 108 13.0037
r186 103 126 0.128424
r187 103 105 6.16843
r188 102 125 0.494161
r189 101 127 0.494161
r190 101 102 4.58464
r191 99 139 1.16709
r192 97 125 0.128424
r193 97 99 2.16729
r194 95 126 0.494161
r195 95 96 7.46046
r196 93 134 1.16709
r197 91 96 0.652036
r198 91 93 2.16729
r199 87 124 0.306046
r200 87 89 1.82344
r201 85 125 0.494161
r202 85 86 10.1279
r203 84 124 0.349767
r204 83 86 0.652036
r205 83 84 5.50157
r206 81 117 1.16709
r207 77 105 1.16709
r208 72 89 1.16709
r209 64 148 0.0476429
r210 64 66 1.92555
r211 59 66 0.5835
r212 58 60 0.652036
r213 58 59 2.8008
r214 55 66 0.0685365
r215 51 139 0.0476429
r216 49 51 1.45875
r217 48 52 0.652036
r218 48 51 1.45875
r219 45 49 0.652036
r220 41 134 0.0476429
r221 39 41 1.45875
r222 38 42 0.652036
r223 38 41 1.45875
r224 35 39 0.652036
r225 20 81 0.123773
r226 18 60 5.1348
r227 16 77 0.123773
r228 14 55 5.1348
r229 12 77 0.123773
r230 10 52 5.1348
r231 8 45 5.1348
r232 6 35 5.1348
r233 4 42 5.1348
r234 2 72 0.123773
.ends

.subckt PM_G4_MUX2_N3_VSS 2 4 6 8 10 12 14 16 18 20 38 39 41 48 49 59 72 77 81
+ 84 89 94 99 104 109 118 123 132 140 141 146 152 153 158 164 170 172 177 179
+ 181 182 183 184 185 Vss
c124 185 Vss 4.28045e-19
c125 184 Vss 3.62111e-19
c126 183 Vss 3.91906e-19
c127 182 Vss 3.21876e-19
c128 179 Vss 0.00582395f
c129 177 Vss 0.00193102f
c130 172 Vss 0.00135159f
c131 170 Vss 0.00259462f
c132 164 Vss 0.00592925f
c133 158 Vss 0.00385718f
c134 153 Vss 5.94991e-19
c135 152 Vss 0.00258264f
c136 147 Vss 0.00135554f
c137 146 Vss 0.00523922f
c138 141 Vss 0.00344346f
c139 140 Vss 0.00104615f
c140 132 Vss 0.00918942f
c141 123 Vss 0.00383026f
c142 118 Vss 0.00413434f
c143 109 Vss 3.63432e-19
c144 104 Vss 0.0017597f
c145 99 Vss 0.00131312f
c146 94 Vss 6.11605e-19
c147 89 Vss 0.00100326f
c148 84 Vss 0.00146588f
c149 81 Vss 0.00807726f
c150 77 Vss 0.00622224f
c151 72 Vss 0.0101685f
c152 65 Vss 0.0783825f
c153 59 Vss 0.0350566f
c154 58 Vss 0.0688416f
c155 49 Vss 0.0347733f
c156 48 Vss 0.100364f
c157 41 Vss 8.95828e-20
c158 39 Vss 0.0350852f
c159 38 Vss 0.0994129f
c160 20 Vss 0.190105f
c161 16 Vss 0.189529f
c162 14 Vss 0.00143493f
c163 12 Vss 0.189243f
c164 10 Vss 0.189689f
c165 4 Vss 0.190073f
c166 2 Vss 0.189016f
r167 178 185 0.551426
r168 178 179 18.3386
r169 177 185 0.551426
r170 176 177 5.50157
r171 172 185 0.0828784
r172 171 184 0.494161
r173 170 179 0.652036
r174 170 171 4.41793
r175 166 184 0.128424
r176 165 183 0.494161
r177 164 176 0.652036
r178 164 165 13.0037
r179 160 183 0.128424
r180 159 182 0.494161
r181 158 184 0.494161
r182 158 159 10.2946
r183 154 182 0.128424
r184 152 183 0.494161
r185 152 153 7.46046
r186 148 153 0.652036
r187 146 182 0.494161
r188 146 147 10.1279
r189 142 181 0.306046
r190 141 147 0.652036
r191 140 181 0.349767
r192 140 141 5.50157
r193 109 172 1.82344
r194 104 132 1.16709
r195 104 166 2.16729
r196 99 160 6.16843
r197 94 123 1.16709
r198 94 154 2.16729
r199 89 118 1.16709
r200 89 148 2.16729
r201 84 142 1.82344
r202 81 109 1.16709
r203 77 99 1.16709
r204 72 84 1.16709
r205 65 132 0.0476429
r206 63 65 1.8672
r207 60 63 0.0685365
r208 58 63 0.5835
r209 58 59 2.8008
r210 55 59 0.652036
r211 51 123 0.0476429
r212 49 51 1.45875
r213 48 52 0.652036
r214 48 51 1.45875
r215 45 49 0.652036
r216 41 118 0.0476429
r217 39 41 1.45875
r218 38 42 0.652036
r219 38 41 1.45875
r220 35 39 0.652036
r221 20 60 5.1348
r222 18 81 0.123773
r223 16 55 5.1348
r224 14 77 0.123773
r225 12 52 5.1348
r226 10 45 5.1348
r227 8 77 0.123773
r228 6 72 0.123773
r229 4 35 5.1348
r230 2 42 5.1348
.ends

.subckt PM_G4_MUX2_N3_ZI 2 4 6 8 10 12 27 28 43 47 50 55 60 65 81 82 91 Vss
c65 82 Vss 9.82283e-19
c66 81 Vss 0.00344769f
c67 65 Vss 0.00531208f
c68 60 Vss 0.00107621f
c69 55 Vss 0.00120586f
c70 50 Vss 0.00184713f
c71 47 Vss 0.00665316f
c72 43 Vss 0.00665316f
c73 28 Vss 0.206957f
c74 27 Vss 8.47557e-20
c75 23 Vss 0.0247918f
c76 12 Vss 0.00143493f
c77 10 Vss 0.00143493f
c78 4 Vss 0.189507f
c79 2 Vss 0.180667f
r80 87 91 0.494161
r81 83 91 0.494161
r82 81 91 0.128424
r83 81 82 13.2121
r84 77 82 0.652036
r85 60 87 5.50157
r86 55 83 6.16843
r87 50 65 1.16709
r88 50 77 2.16729
r89 47 60 1.16709
r90 43 55 1.16709
r91 31 65 0.0476429
r92 29 31 0.326018
r93 29 31 0.1167
r94 28 32 0.652036
r95 28 31 6.7686
r96 27 65 0.357321
r97 23 31 0.326018
r98 23 27 0.40845
r99 12 47 0.123773
r100 10 43 0.123773
r101 8 47 0.123773
r102 6 43 0.123773
r103 4 32 5.1348
r104 2 27 4.72635
.ends

.subckt PM_G4_MUX2_N3_Z 2 4 13 16 Vss
c13 16 Vss 2.03714e-19
c14 13 Vss 0.00452755f
c15 4 Vss 0.00143493f
r16 16 19 0.0416786
r17 13 19 1.16709
r18 4 13 0.123773
r19 2 13 0.123773
.ends

.subckt PM_G4_MUX2_N3_SELI 2 4 6 8 18 21 29 33 36 38 43 44 52 57 71 76 77 Vss
c72 77 Vss 8.29462e-19
c73 76 Vss 1.71087e-19
c74 71 Vss 0.00163664f
c75 57 Vss 0.00292618f
c76 52 Vss 0.00318194f
c77 44 Vss 0.00264419f
c78 43 Vss 8.75265e-19
c79 38 Vss 0.00210957f
c80 36 Vss 3.78531e-19
c81 33 Vss 0.00302148f
c82 29 Vss 0.00524134f
c83 21 Vss 0.16662f
c84 18 Vss 7.81442e-20
c85 6 Vss 0.166657f
c86 4 Vss 0.00143493f
r87 76 77 0.655813
r88 75 76 3.501
r89 71 75 0.655813
r90 43 52 1.16709
r91 43 71 2.00578
r92 43 44 0.513084
r93 38 57 1.16709
r94 38 77 2.00578
r95 36 44 7.46046
r96 31 36 0.652036
r97 31 33 7.91893
r98 29 33 1.16709
r99 21 57 0.50025
r100 18 52 0.50025
r101 8 21 4.37625
r102 6 18 4.37625
r103 4 29 0.123773
r104 2 29 0.123773
.ends

.subckt PM_G4_MUX2_N3_SEL 2 4 6 8 16 17 22 26 33 36 40 41 44 45 47 49 56 57 59
+ 64 69 Vss
c65 69 Vss 0.00293892f
c66 64 Vss 0.00330355f
c67 59 Vss 0.00281287f
c68 57 Vss 3.29949e-19
c69 56 Vss 0.00195862f
c70 49 Vss 4.84367e-19
c71 47 Vss 0.00164668f
c72 45 Vss 5.48919e-19
c73 44 Vss 0.00192809f
c74 41 Vss 0.00187197f
c75 36 Vss 8.44333e-20
c76 33 Vss 9.14819e-20
c77 26 Vss 0.16662f
c78 22 Vss 0.180313f
c79 20 Vss 0.0247918f
c80 17 Vss 0.0358843f
c81 16 Vss 0.179072f
c82 8 Vss 0.16662f
c83 2 Vss 0.193774f
r84 55 64 1.16709
r85 55 57 0.4602
r86 55 56 0.52504
r87 52 59 1.16709
r88 49 52 0.5835
r89 47 69 1.16709
r90 45 47 2.00578
r91 43 45 0.655813
r92 43 44 3.501
r93 41 44 0.655813
r94 41 57 1.49522
r95 40 56 2.58407
r96 38 49 0.0685365
r97 38 40 2.00057
r98 36 59 0.0476429
r99 33 69 0.50025
r100 26 64 0.50025
r101 22 59 0.357321
r102 20 36 0.326018
r103 20 22 0.40845
r104 17 36 6.7686
r105 16 36 0.326018
r106 16 36 0.1167
r107 13 17 0.652036
r108 8 33 4.37625
r109 6 26 4.37625
r110 4 22 4.72635
r111 2 13 5.1348
.ends

.subckt PM_G4_MUX2_N3_B 2 4 14 17 20 23 Vss
c30 23 Vss 0.00439028f
c31 20 Vss 2.87096e-19
c32 14 Vss 0.0853197f
c33 2 Vss 0.656289f
r34 20 23 1.16709
r35 17 20 0.109406
r36 14 23 0.0476429
r37 11 14 1.92555
r38 7 11 0.0685365
r39 4 7 5.1348
r40 2 4 17.9718
.ends

.subckt PM_G4_MUX2_N3_A 2 4 12 14 20 23 Vss
c24 23 Vss 0.00548676f
c25 20 Vss 2.95003e-19
c26 14 Vss 0.0835366f
c27 12 Vss 8.63834e-20
c28 2 Vss 0.664171f
r29 17 23 1.16709
r30 17 20 0.0364688
r31 12 23 0.0476429
r32 12 14 1.92555
r33 7 14 0.0685365
r34 2 4 17.9718
r35 2 7 5.1348
.ends

.subckt G4_MUX2_N3  VDD VSS Z SEL B A
*
* A	A
* B	B
* SEL	SEL
* Z	Z
* VSS	VSS
* VDD	VDD
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_ZI_XI6.X0_CG N_VSS_XI6.X0_PGS
+ N_VDD_XI6.X0_S TIGFET_HPNW12
XI12.X0 N_SELI_XI12.X0_D N_VDD_XI12.X0_PGD N_SEL_XI12.X0_CG N_VDD_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW12
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_ZI_XI5.X0_CG N_VDD_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW12
XI13.X0 N_SELI_XI13.X0_D N_VSS_XI13.X0_PGD N_SEL_XI13.X0_CG N_VSS_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW12
XI17.X0 N_ZI_XI17.X0_D N_VDD_XI17.X0_PGD N_SELI_XI17.X0_CG N_B_XI17.X0_PGS
+ N_VSS_XI17.X0_S TIGFET_HPNW12
XI15.X0 N_ZI_XI15.X0_D N_VSS_XI15.X0_PGD N_SEL_XI15.X0_CG N_B_XI15.X0_PGS
+ N_VDD_XI15.X0_S TIGFET_HPNW12
XI16.X0 N_ZI_XI16.X0_D N_VDD_XI16.X0_PGD N_SEL_XI16.X0_CG N_A_XI16.X0_PGS
+ N_VSS_XI16.X0_S TIGFET_HPNW12
XI14.X0 N_ZI_XI14.X0_D N_VSS_XI14.X0_PGD N_SELI_XI14.X0_CG N_A_XI14.X0_PGS
+ N_VDD_XI14.X0_S TIGFET_HPNW12
*
x_PM_G4_MUX2_N3_VDD N_VDD_XI6.X0_S N_VDD_XI12.X0_PGD N_VDD_XI12.X0_PGS
+ N_VDD_XI5.X0_PGD N_VDD_XI5.X0_PGS N_VDD_XI13.X0_S N_VDD_XI17.X0_PGD
+ N_VDD_XI15.X0_S N_VDD_XI16.X0_PGD N_VDD_XI14.X0_S N_VDD_c_12_p N_VDD_c_8_p
+ N_VDD_c_102_p N_VDD_c_127_p N_VDD_c_92_p N_VDD_c_86_p N_VDD_c_15_p
+ N_VDD_c_74_p N_VDD_c_10_p N_VDD_c_9_p N_VDD_c_17_p N_VDD_c_22_p N_VDD_c_13_p
+ N_VDD_c_49_p N_VDD_c_20_p N_VDD_c_16_p N_VDD_c_5_p N_VDD_c_14_p N_VDD_c_29_p
+ N_VDD_c_34_p N_VDD_c_61_p N_VDD_c_30_p N_VDD_c_33_p VDD N_VDD_c_52_p
+ N_VDD_c_56_p N_VDD_c_59_p N_VDD_c_66_p N_VDD_c_25_p N_VDD_c_21_p N_VDD_c_100_p
+ Vss PM_G4_MUX2_N3_VDD
x_PM_G4_MUX2_N3_VSS N_VSS_XI6.X0_PGD N_VSS_XI6.X0_PGS N_VSS_XI12.X0_S
+ N_VSS_XI5.X0_S N_VSS_XI13.X0_PGD N_VSS_XI13.X0_PGS N_VSS_XI17.X0_S
+ N_VSS_XI15.X0_PGD N_VSS_XI16.X0_S N_VSS_XI14.X0_PGD N_VSS_c_139_n
+ N_VSS_c_141_n N_VSS_c_202_p N_VSS_c_246_p N_VSS_c_143_n N_VSS_c_145_n
+ N_VSS_c_226_p N_VSS_c_146_n N_VSS_c_205_p N_VSS_c_148_n N_VSS_c_149_n
+ N_VSS_c_153_n N_VSS_c_157_n N_VSS_c_162_n N_VSS_c_165_n N_VSS_c_167_n
+ N_VSS_c_170_n N_VSS_c_174_n N_VSS_c_176_n N_VSS_c_177_n N_VSS_c_179_n
+ N_VSS_c_181_n N_VSS_c_184_n N_VSS_c_185_n N_VSS_c_188_n N_VSS_c_191_n
+ N_VSS_c_192_n N_VSS_c_193_n N_VSS_c_194_n VSS N_VSS_c_198_n N_VSS_c_199_n
+ N_VSS_c_200_n N_VSS_c_201_n Vss PM_G4_MUX2_N3_VSS
x_PM_G4_MUX2_N3_ZI N_ZI_XI6.X0_CG N_ZI_XI5.X0_CG N_ZI_XI17.X0_D N_ZI_XI15.X0_D
+ N_ZI_XI16.X0_D N_ZI_XI14.X0_D N_ZI_c_271_n N_ZI_c_256_n N_ZI_c_257_n
+ N_ZI_c_258_n N_ZI_c_276_n N_ZI_c_262_n N_ZI_c_264_n N_ZI_c_296_p N_ZI_c_270_n
+ N_ZI_c_290_n N_ZI_c_306_p Vss PM_G4_MUX2_N3_ZI
x_PM_G4_MUX2_N3_Z N_Z_XI6.X0_D N_Z_XI5.X0_D N_Z_c_321_n Z Vss PM_G4_MUX2_N3_Z
x_PM_G4_MUX2_N3_SELI N_SELI_XI12.X0_D N_SELI_XI13.X0_D N_SELI_XI17.X0_CG
+ N_SELI_XI14.X0_CG N_SELI_c_334_n N_SELI_c_404_p N_SELI_c_335_n N_SELI_c_338_n
+ N_SELI_c_361_n N_SELI_c_341_n N_SELI_c_342_n N_SELI_c_343_n N_SELI_c_346_n
+ N_SELI_c_347_n N_SELI_c_357_n N_SELI_c_371_n N_SELI_c_374_n Vss
+ PM_G4_MUX2_N3_SELI
x_PM_G4_MUX2_N3_SEL N_SEL_XI12.X0_CG N_SEL_XI13.X0_CG N_SEL_XI15.X0_CG
+ N_SEL_XI16.X0_CG N_SEL_c_406_n N_SEL_c_422_n N_SEL_c_456_p N_SEL_c_457_p
+ N_SEL_c_467_p N_SEL_c_415_n SEL N_SEL_c_407_n N_SEL_c_408_n N_SEL_c_429_n
+ N_SEL_c_409_n N_SEL_c_418_n N_SEL_c_411_n N_SEL_c_445_n N_SEL_c_420_n
+ N_SEL_c_448_n N_SEL_c_413_n Vss PM_G4_MUX2_N3_SEL
x_PM_G4_MUX2_N3_B N_B_XI17.X0_PGS N_B_XI15.X0_PGS N_B_c_477_n B N_B_c_471_n
+ N_B_c_473_n Vss PM_G4_MUX2_N3_B
x_PM_G4_MUX2_N3_A N_A_XI16.X0_PGS N_A_XI14.X0_PGS N_A_c_520_n N_A_c_503_n A
+ N_A_c_509_n Vss PM_G4_MUX2_N3_A
cc_1 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.00200866f
cc_2 N_VDD_XI12.X0_PGS N_VSS_XI6.X0_PGS 2.44446e-19
cc_3 N_VDD_XI12.X0_PGD N_VSS_XI13.X0_PGD 0.00195824f
cc_4 N_VDD_XI5.X0_PGS N_VSS_XI13.X0_PGS 2.27381e-19
cc_5 N_VDD_c_5_p N_VSS_XI13.X0_PGS 2.10824e-19
cc_6 N_VDD_XI17.X0_PGD N_VSS_XI15.X0_PGD 2.31533e-19
cc_7 N_VDD_XI16.X0_PGD N_VSS_XI14.X0_PGD 2.31533e-19
cc_8 N_VDD_c_8_p N_VSS_c_139_n 0.00200866f
cc_9 N_VDD_c_9_p N_VSS_c_139_n 3.89167e-19
cc_10 N_VDD_c_10_p N_VSS_c_141_n 4.28478e-19
cc_11 N_VDD_c_9_p N_VSS_c_141_n 4.0633e-19
cc_12 N_VDD_c_12_p N_VSS_c_143_n 0.00195824f
cc_13 N_VDD_c_13_p N_VSS_c_143_n 3.10186e-19
cc_14 N_VDD_c_14_p N_VSS_c_145_n 9.06483e-19
cc_15 N_VDD_c_15_p N_VSS_c_146_n 3.23931e-19
cc_16 N_VDD_c_16_p N_VSS_c_146_n 2.74986e-19
cc_17 N_VDD_c_17_p N_VSS_c_148_n 4.89302e-19
cc_18 N_VDD_c_10_p N_VSS_c_149_n 8.67538e-19
cc_19 N_VDD_c_9_p N_VSS_c_149_n 0.00141228f
cc_20 N_VDD_c_20_p N_VSS_c_149_n 8.83788e-19
cc_21 N_VDD_c_21_p N_VSS_c_149_n 3.48267e-19
cc_22 N_VDD_c_22_p N_VSS_c_153_n 8.50587e-19
cc_23 N_VDD_c_13_p N_VSS_c_153_n 0.00141228f
cc_24 N_VDD_c_5_p N_VSS_c_153_n 0.00180638f
cc_25 N_VDD_c_25_p N_VSS_c_153_n 3.48267e-19
cc_26 N_VDD_c_10_p N_VSS_c_157_n 2.85826e-19
cc_27 N_VDD_c_20_p N_VSS_c_157_n 3.92901e-19
cc_28 N_VDD_c_16_p N_VSS_c_157_n 2.9533e-19
cc_29 N_VDD_c_29_p N_VSS_c_157_n 7.06793e-19
cc_30 N_VDD_c_30_p N_VSS_c_157_n 4.71075e-19
cc_31 N_VDD_c_5_p N_VSS_c_162_n 2.93442e-19
cc_32 N_VDD_c_14_p N_VSS_c_162_n 0.00161703f
cc_33 N_VDD_c_33_p N_VSS_c_162_n 4.28751e-19
cc_34 N_VDD_c_34_p N_VSS_c_165_n 3.5277e-19
cc_35 N_VDD_c_30_p N_VSS_c_165_n 0.00187494f
cc_36 N_VDD_c_10_p N_VSS_c_167_n 3.66936e-19
cc_37 N_VDD_c_9_p N_VSS_c_167_n 0.00114511f
cc_38 N_VDD_c_21_p N_VSS_c_167_n 6.489e-19
cc_39 N_VDD_c_22_p N_VSS_c_170_n 3.82294e-19
cc_40 N_VDD_c_13_p N_VSS_c_170_n 0.00114511f
cc_41 N_VDD_c_5_p N_VSS_c_170_n 9.55349e-19
cc_42 N_VDD_c_25_p N_VSS_c_170_n 6.46219e-19
cc_43 N_VDD_c_14_p N_VSS_c_174_n 2.26455e-19
cc_44 N_VDD_c_33_p N_VSS_c_174_n 5.86293e-19
cc_45 N_VDD_c_10_p N_VSS_c_176_n 3.30364e-19
cc_46 N_VDD_c_22_p N_VSS_c_177_n 3.85245e-19
cc_47 N_VDD_c_5_p N_VSS_c_177_n 2.91233e-19
cc_48 N_VDD_c_13_p N_VSS_c_179_n 0.00427835f
cc_49 N_VDD_c_49_p N_VSS_c_179_n 0.00166784f
cc_50 N_VDD_c_9_p N_VSS_c_181_n 0.00425881f
cc_51 N_VDD_c_16_p N_VSS_c_181_n 0.00135965f
cc_52 N_VDD_c_52_p N_VSS_c_181_n 0.0010575f
cc_53 N_VDD_c_9_p N_VSS_c_184_n 0.00176255f
cc_54 N_VDD_c_13_p N_VSS_c_185_n 0.00138037f
cc_55 N_VDD_c_14_p N_VSS_c_185_n 0.00614137f
cc_56 N_VDD_c_56_p N_VSS_c_185_n 0.00120833f
cc_57 N_VDD_c_16_p N_VSS_c_188_n 0.00135965f
cc_58 N_VDD_c_34_p N_VSS_c_188_n 0.00823017f
cc_59 N_VDD_c_59_p N_VSS_c_188_n 0.00103007f
cc_60 N_VDD_c_14_p N_VSS_c_191_n 0.00457914f
cc_61 N_VDD_c_61_p N_VSS_c_192_n 4.01154e-19
cc_62 N_VDD_c_30_p N_VSS_c_193_n 0.0041789f
cc_63 N_VDD_c_5_p N_VSS_c_194_n 4.46614e-19
cc_64 N_VDD_c_30_p N_VSS_c_194_n 0.00867926f
cc_65 N_VDD_c_33_p N_VSS_c_194_n 0.00355235f
cc_66 N_VDD_c_66_p N_VSS_c_194_n 0.0010706f
cc_67 N_VDD_c_13_p N_VSS_c_198_n 7.23159e-19
cc_68 N_VDD_c_16_p N_VSS_c_199_n 0.00111918f
cc_69 N_VDD_c_14_p N_VSS_c_200_n 7.61747e-19
cc_70 N_VDD_c_30_p N_VSS_c_201_n 9.16632e-19
cc_71 N_VDD_XI5.X0_PGD N_ZI_c_256_n 3.96029e-19
cc_72 N_VDD_c_34_p N_ZI_c_257_n 2.74986e-19
cc_73 N_VDD_c_15_p N_ZI_c_258_n 3.43419e-19
cc_74 N_VDD_c_74_p N_ZI_c_258_n 3.43419e-19
cc_75 N_VDD_c_5_p N_ZI_c_258_n 3.48267e-19
cc_76 N_VDD_c_61_p N_ZI_c_258_n 3.72199e-19
cc_77 N_VDD_c_34_p N_ZI_c_262_n 2.9533e-19
cc_78 N_VDD_c_30_p N_ZI_c_262_n 9.20678e-19
cc_79 N_VDD_c_15_p N_ZI_c_264_n 3.48267e-19
cc_80 N_VDD_c_74_p N_ZI_c_264_n 3.48267e-19
cc_81 N_VDD_c_5_p N_ZI_c_264_n 4.99861e-19
cc_82 N_VDD_c_14_p N_ZI_c_264_n 3.21336e-19
cc_83 N_VDD_c_61_p N_ZI_c_264_n 5.226e-19
cc_84 N_VDD_c_30_p N_ZI_c_264_n 2.34601e-19
cc_85 N_VDD_c_13_p N_ZI_c_270_n 2.91231e-19
cc_86 N_VDD_c_86_p N_Z_c_321_n 3.43419e-19
cc_87 N_VDD_c_9_p N_Z_c_321_n 2.74986e-19
cc_88 N_VDD_c_17_p N_Z_c_321_n 3.72199e-19
cc_89 N_VDD_c_86_p Z 3.48267e-19
cc_90 N_VDD_c_9_p Z 3.66281e-19
cc_91 N_VDD_c_17_p Z 7.4527e-19
cc_92 N_VDD_c_92_p N_SELI_c_334_n 4.99294e-19
cc_93 N_VDD_c_15_p N_SELI_c_335_n 3.43419e-19
cc_94 N_VDD_c_13_p N_SELI_c_335_n 2.74986e-19
cc_95 N_VDD_c_5_p N_SELI_c_335_n 3.48267e-19
cc_96 N_VDD_c_15_p N_SELI_c_338_n 3.48267e-19
cc_97 N_VDD_c_13_p N_SELI_c_338_n 3.8357e-19
cc_98 N_VDD_c_5_p N_SELI_c_338_n 6.94315e-19
cc_99 N_VDD_c_30_p N_SELI_c_341_n 4.32468e-19
cc_100 N_VDD_c_100_p N_SELI_c_342_n 2.17157e-19
cc_101 N_VDD_XI5.X0_PGD N_SELI_c_343_n 2.35597e-19
cc_102 N_VDD_c_102_p N_SELI_c_343_n 2.28823e-19
cc_103 N_VDD_c_20_p N_SELI_c_343_n 2.91405e-19
cc_104 N_VDD_c_29_p N_SELI_c_346_n 2.28697e-19
cc_105 N_VDD_c_30_p N_SELI_c_347_n 3.66936e-19
cc_106 N_VDD_XI12.X0_PGD N_SEL_c_406_n 4.09718e-19
cc_107 N_VDD_c_14_p N_SEL_c_407_n 3.4535e-19
cc_108 N_VDD_c_30_p N_SEL_c_408_n 5.4414e-19
cc_109 N_VDD_c_34_p N_SEL_c_409_n 3.57377e-19
cc_110 N_VDD_c_30_p N_SEL_c_409_n 5.05119e-19
cc_111 N_VDD_c_15_p N_SEL_c_411_n 4.75243e-19
cc_112 N_VDD_c_5_p N_SEL_c_411_n 7.80048e-19
cc_113 N_VDD_c_30_p N_SEL_c_413_n 3.66936e-19
cc_114 N_VDD_c_5_p N_B_c_471_n 0.00142218f
cc_115 N_VDD_c_14_p N_B_c_471_n 0.00141439f
cc_116 N_VDD_c_5_p N_B_c_473_n 9.67317e-19
cc_117 N_VDD_c_14_p N_B_c_473_n 0.00120343f
cc_118 N_VDD_XI16.X0_PGD N_A_XI16.X0_PGS 0.00146246f
cc_119 N_VDD_c_30_p N_A_XI16.X0_PGS 0.00124298f
cc_120 N_VDD_c_34_p N_A_c_503_n 3.5103e-19
cc_121 N_VDD_c_30_p N_A_c_503_n 3.92527e-19
cc_122 N_VDD_c_29_p A 5.27373e-19
cc_123 N_VDD_c_34_p A 0.00141439f
cc_124 N_VDD_c_30_p A 5.12828e-19
cc_125 N_VDD_c_100_p A 3.44698e-19
cc_126 N_VDD_XI16.X0_PGD N_A_c_509_n 3.32271e-19
cc_127 N_VDD_c_127_p N_A_c_509_n 0.00480616f
cc_128 N_VDD_c_29_p N_A_c_509_n 3.95721e-19
cc_129 N_VDD_c_34_p N_A_c_509_n 0.00120343f
cc_130 N_VDD_c_30_p N_A_c_509_n 3.70842e-19
cc_131 N_VDD_c_100_p N_A_c_509_n 6.02643e-19
cc_132 N_VSS_c_202_p N_ZI_c_271_n 5.35095e-19
cc_133 N_VSS_XI6.X0_PGD N_ZI_c_256_n 4.09718e-19
cc_134 N_VSS_c_146_n N_ZI_c_257_n 3.43419e-19
cc_135 N_VSS_c_205_p N_ZI_c_257_n 3.43419e-19
cc_136 N_VSS_c_165_n N_ZI_c_257_n 3.48267e-19
cc_137 N_VSS_c_149_n N_ZI_c_276_n 3.27284e-19
cc_138 N_VSS_c_167_n N_ZI_c_276_n 2.15082e-19
cc_139 N_VSS_c_146_n N_ZI_c_262_n 3.48267e-19
cc_140 N_VSS_c_205_p N_ZI_c_262_n 3.48267e-19
cc_141 N_VSS_c_157_n N_ZI_c_262_n 0.00100597f
cc_142 N_VSS_c_165_n N_ZI_c_262_n 4.40384e-19
cc_143 N_VSS_c_188_n N_ZI_c_262_n 3.80707e-19
cc_144 N_VSS_c_192_n N_ZI_c_262_n 6.1924e-19
cc_145 N_VSS_c_194_n N_ZI_c_262_n 0.00228731f
cc_146 N_VSS_c_185_n N_ZI_c_264_n 3.80707e-19
cc_147 N_VSS_c_153_n N_ZI_c_270_n 2.70732e-19
cc_148 N_VSS_c_157_n N_ZI_c_270_n 4.41808e-19
cc_149 N_VSS_c_181_n N_ZI_c_270_n 7.14893e-19
cc_150 N_VSS_c_185_n N_ZI_c_270_n 0.00105381f
cc_151 N_VSS_c_179_n N_ZI_c_290_n 7.92312e-19
cc_152 N_VSS_c_146_n N_Z_c_321_n 3.43419e-19
cc_153 N_VSS_c_157_n N_Z_c_321_n 3.48267e-19
cc_154 N_VSS_c_146_n Z 3.48267e-19
cc_155 N_VSS_c_157_n Z 7.85754e-19
cc_156 N_VSS_c_226_p N_SELI_c_335_n 3.43419e-19
cc_157 N_VSS_c_148_n N_SELI_c_335_n 3.48267e-19
cc_158 N_VSS_c_226_p N_SELI_c_338_n 3.48267e-19
cc_159 N_VSS_c_148_n N_SELI_c_338_n 5.71987e-19
cc_160 N_VSS_c_194_n N_SELI_c_341_n 6.69121e-19
cc_161 N_VSS_c_146_n N_SELI_c_343_n 5.11666e-19
cc_162 N_VSS_c_157_n N_SELI_c_343_n 6.75781e-19
cc_163 N_VSS_c_181_n N_SELI_c_343_n 3.61249e-19
cc_164 N_VSS_c_174_n N_SELI_c_347_n 5.05931e-19
cc_165 N_VSS_c_188_n N_SELI_c_357_n 6.42552e-19
cc_166 N_VSS_c_194_n N_SELI_c_357_n 6.85767e-19
cc_167 N_VSS_XI13.X0_PGD N_SEL_c_406_n 4.03539e-19
cc_168 N_VSS_c_170_n N_SEL_c_415_n 5.28949e-19
cc_169 N_VSS_c_194_n N_SEL_c_408_n 2.60801e-19
cc_170 N_VSS_c_188_n N_SEL_c_409_n 2.29905e-19
cc_171 N_VSS_c_170_n N_SEL_c_418_n 2.18943e-19
cc_172 N_VSS_c_185_n N_SEL_c_411_n 3.31177e-19
cc_173 N_VSS_c_153_n N_SEL_c_420_n 2.15082e-19
cc_174 N_VSS_XI13.X0_PGS N_B_XI17.X0_PGS 0.00187616f
cc_175 N_VSS_XI15.X0_PGD N_B_XI17.X0_PGS 0.00145666f
cc_176 N_VSS_c_246_p N_B_c_477_n 0.00187616f
cc_177 N_VSS_c_162_n N_B_c_471_n 3.92469e-19
cc_178 N_VSS_c_174_n N_B_c_471_n 3.5189e-19
cc_179 N_VSS_c_185_n N_B_c_471_n 2.15119e-19
cc_180 N_VSS_XI15.X0_PGD N_B_c_473_n 3.23173e-19
cc_181 N_VSS_c_145_n N_B_c_473_n 0.00295829f
cc_182 N_VSS_c_162_n N_B_c_473_n 3.5189e-19
cc_183 N_VSS_c_170_n N_B_c_473_n 6.40394e-19
cc_184 N_VSS_c_174_n N_B_c_473_n 6.81736e-19
cc_185 N_VSS_c_188_n A 2.41977e-19
cc_186 N_ZI_c_256_n N_Z_c_321_n 6.90199e-19
cc_187 N_ZI_c_264_n N_SELI_c_338_n 9.22717e-19
cc_188 N_ZI_c_270_n N_SELI_c_338_n 0.00230161f
cc_189 N_ZI_c_256_n N_SELI_c_361_n 3.69647e-19
cc_190 N_ZI_c_276_n N_SELI_c_361_n 0.00194838f
cc_191 N_ZI_c_296_p N_SELI_c_361_n 9.76295e-19
cc_192 N_ZI_c_264_n N_SELI_c_341_n 0.00164769f
cc_193 N_ZI_c_262_n N_SELI_c_342_n 0.00166362f
cc_194 N_ZI_c_270_n N_SELI_c_342_n 0.00145462f
cc_195 N_ZI_c_256_n N_SELI_c_343_n 8.08917e-19
cc_196 N_ZI_c_270_n N_SELI_c_343_n 0.0018158f
cc_197 N_ZI_c_262_n N_SELI_c_357_n 7.72596e-19
cc_198 N_ZI_c_270_n N_SELI_c_357_n 7.93892e-19
cc_199 N_ZI_c_262_n N_SELI_c_371_n 6.01706e-19
cc_200 N_ZI_c_264_n N_SELI_c_371_n 3.05282e-19
cc_201 N_ZI_c_306_p N_SELI_c_371_n 6.45182e-19
cc_202 N_ZI_c_264_n N_SELI_c_374_n 8.28497e-19
cc_203 N_ZI_c_256_n N_SEL_c_406_n 0.0037589f
cc_204 N_ZI_c_296_p N_SEL_c_422_n 5.93636e-19
cc_205 N_ZI_c_258_n N_SEL_c_407_n 6.40197e-19
cc_206 N_ZI_c_264_n N_SEL_c_407_n 0.00209308f
cc_207 N_ZI_c_270_n N_SEL_c_407_n 8.88094e-19
cc_208 N_ZI_c_262_n N_SEL_c_408_n 9.51454e-19
cc_209 N_ZI_c_264_n N_SEL_c_408_n 4.59089e-19
cc_210 N_ZI_c_306_p N_SEL_c_408_n 0.00107464f
cc_211 N_ZI_c_257_n N_SEL_c_429_n 6.40197e-19
cc_212 N_ZI_c_262_n N_SEL_c_429_n 0.00193202f
cc_213 N_ZI_c_270_n N_SEL_c_418_n 0.0016105f
cc_214 N_ZI_c_256_n N_SEL_c_420_n 0.00117386f
cc_215 N_ZI_XI5.X0_CG N_B_XI17.X0_PGS 0.0018458f
cc_216 N_Z_c_321_n N_SELI_c_361_n 5.76103e-19
cc_217 Z N_SELI_c_361_n 8.85628e-19
cc_218 N_SELI_c_335_n N_SEL_c_406_n 6.90199e-19
cc_219 N_SELI_c_338_n N_SEL_c_406_n 8.57466e-19
cc_220 N_SELI_c_343_n N_SEL_c_406_n 2.79929e-19
cc_221 N_SELI_c_341_n N_SEL_c_407_n 0.00141479f
cc_222 N_SELI_c_347_n N_SEL_c_407_n 9.76295e-19
cc_223 N_SELI_c_338_n N_SEL_c_408_n 3.66824e-19
cc_224 N_SELI_c_342_n N_SEL_c_429_n 0.00170409f
cc_225 N_SELI_c_346_n N_SEL_c_429_n 9.29204e-19
cc_226 N_SELI_c_341_n N_SEL_c_409_n 9.15421e-19
cc_227 N_SELI_c_338_n N_SEL_c_418_n 0.00216212f
cc_228 N_SELI_c_343_n N_SEL_c_418_n 7.61998e-19
cc_229 N_SELI_c_343_n N_SEL_c_411_n 0.00193122f
cc_230 N_SELI_c_342_n N_SEL_c_445_n 0.00200661f
cc_231 N_SELI_c_338_n N_SEL_c_420_n 0.00109331f
cc_232 N_SELI_c_343_n N_SEL_c_420_n 4.73568e-19
cc_233 N_SELI_c_341_n N_SEL_c_448_n 3.48267e-19
cc_234 N_SELI_c_342_n N_SEL_c_448_n 4.95293e-19
cc_235 N_SELI_c_346_n N_SEL_c_448_n 0.00480115f
cc_236 N_SELI_c_347_n N_SEL_c_448_n 9.11855e-19
cc_237 N_SELI_c_341_n N_SEL_c_413_n 4.56568e-19
cc_238 N_SELI_c_342_n N_SEL_c_413_n 3.48267e-19
cc_239 N_SELI_c_346_n N_SEL_c_413_n 9.03632e-19
cc_240 N_SELI_c_347_n N_SEL_c_413_n 0.00245376f
cc_241 N_SELI_XI17.X0_CG N_B_XI17.X0_PGS 4.83278e-19
cc_242 N_SELI_c_338_n N_B_XI17.X0_PGS 2.54355e-19
cc_243 N_SELI_c_343_n N_B_XI17.X0_PGS 8.44835e-19
cc_244 N_SELI_c_346_n N_B_XI17.X0_PGS 0.00126314f
cc_245 N_SELI_c_404_p N_A_XI16.X0_PGS 4.99479e-19
cc_246 N_SELI_c_347_n N_A_XI16.X0_PGS 0.001089f
cc_247 N_SEL_c_456_p N_B_XI17.X0_PGS 2.07014e-19
cc_248 N_SEL_c_457_p N_B_XI17.X0_PGS 4.77845e-19
cc_249 N_SEL_c_411_n N_B_XI17.X0_PGS 7.43585e-19
cc_250 N_SEL_c_420_n N_B_XI17.X0_PGS 0.00100354f
cc_251 N_SEL_c_448_n N_B_XI17.X0_PGS 0.00142122f
cc_252 N_SEL_c_445_n N_B_c_471_n 2.97827e-19
cc_253 N_SEL_c_448_n N_B_c_471_n 2.15082e-19
cc_254 N_SEL_c_445_n N_B_c_473_n 2.18943e-19
cc_255 N_SEL_c_448_n N_B_c_473_n 5.28949e-19
cc_256 N_SEL_XI16.X0_CG N_A_XI16.X0_PGS 4.99479e-19
cc_257 N_SEL_c_413_n N_A_XI16.X0_PGS 0.001089f
cc_258 N_SEL_c_467_p N_A_c_520_n 5.05931e-19
cc_259 N_SEL_c_409_n A 2.92011e-19
cc_260 N_SEL_c_413_n A 2.15082e-19
cc_261 N_SEL_c_409_n N_A_c_509_n 2.15082e-19
cc_262 N_B_XI17.X0_PGS N_A_XI16.X0_PGS 0.00134425f
*
.ends
*
*
.subckt MUX2_HPNW12 A B S0 Y VDD VSS
xgate (VDD VSS Y S0 B A) G4_MUX2_N3
.ends
*
* File: G3_MUXI2_N3.pex.netlist
* Created: Wed Mar  9 15:24:03 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MUXI2_N3_VSS 2 4 6 8 10 12 14 29 39 51 55 60 63 68 73 78 83 92 101
+ 110 115 121 127 133 135 140 142 144 145 146 147 Vss
c77 147 Vss 4.28045e-19
c78 146 Vss 3.62111e-19
c79 145 Vss 3.75522e-19
c80 142 Vss 0.00603414f
c81 140 Vss 0.00196409f
c82 135 Vss 0.00134915f
c83 133 Vss 0.00261859f
c84 128 Vss 0.00128551f
c85 127 Vss 0.00634725f
c86 121 Vss 0.00397667f
c87 115 Vss 0.00552282f
c88 111 Vss 0.00129855f
c89 110 Vss 0.00492065f
c90 101 Vss 0.00967583f
c91 92 Vss 0.00411469f
c92 83 Vss 2.01624e-19
c93 78 Vss 0.0013136f
c94 73 Vss 0.00223792f
c95 68 Vss 4.13309e-19
c96 63 Vss 0.00127305f
c97 60 Vss 0.00806368f
c98 55 Vss 0.00637385f
c99 51 Vss 0.0100822f
c100 45 Vss 0.0783825f
c101 39 Vss 0.0354115f
c102 38 Vss 0.0688416f
c103 29 Vss 0.0347733f
c104 28 Vss 0.101002f
c105 14 Vss 0.189925f
c106 10 Vss 0.190498f
c107 6 Vss 0.190106f
c108 4 Vss 0.189513f
r109 141 147 0.551426
r110 141 142 18.3386
r111 140 147 0.551426
r112 139 140 5.50157
r113 135 147 0.0828784
r114 134 146 0.494161
r115 133 142 0.652036
r116 133 134 4.41793
r117 129 146 0.128424
r118 127 139 0.652036
r119 127 128 13.0037
r120 123 128 0.652036
r121 122 145 0.494161
r122 121 146 0.494161
r123 121 122 10.2946
r124 117 145 0.128424
r125 116 144 0.326018
r126 115 145 0.494161
r127 115 116 10.1279
r128 110 144 0.326018
r129 109 111 0.655813
r130 109 110 5.50157
r131 83 135 1.82344
r132 78 101 1.16709
r133 78 129 2.16729
r134 73 123 6.16843
r135 68 92 1.16709
r136 68 117 2.16729
r137 63 111 1.82344
r138 60 83 1.16709
r139 55 73 1.16709
r140 51 63 1.16709
r141 45 101 0.0476429
r142 43 45 1.8672
r143 40 43 0.0685365
r144 38 43 0.5835
r145 38 39 2.8008
r146 35 39 0.652036
r147 31 92 0.0476429
r148 29 31 1.45875
r149 28 32 0.652036
r150 28 31 1.45875
r151 25 29 0.652036
r152 14 40 5.1348
r153 12 60 0.123773
r154 10 35 5.1348
r155 8 55 0.123773
r156 6 32 5.1348
r157 4 25 5.1348
r158 2 51 0.123773
.ends

.subckt PM_G3_MUXI2_N3_VDD 2 4 6 8 10 12 14 28 38 44 52 56 60 62 63 66 68 72 74
+ 75 76 81 83 84 85 87 89 98 Vss
c91 98 Vss 0.0111734f
c92 89 Vss 0.00463585f
c93 85 Vss 4.52364e-19
c94 84 Vss 4.43941e-19
c95 83 Vss 0.00378478f
c96 81 Vss 0.0102529f
c97 76 Vss 0.00177107f
c98 75 Vss 6.09322e-19
c99 74 Vss 0.0063331f
c100 72 Vss 0.00100496f
c101 68 Vss 0.00791367f
c102 66 Vss 0.00123499f
c103 63 Vss 6.1175e-19
c104 62 Vss 0.00364703f
c105 60 Vss 8.24271e-19
c106 56 Vss 0.00850511f
c107 52 Vss 0.00631561f
c108 39 Vss 0.0806024f
c109 38 Vss 0.103898f
c110 29 Vss 0.0367394f
c111 28 Vss 0.101312f
c112 12 Vss 0.189418f
c113 10 Vss 0.00143493f
c114 8 Vss 0.191033f
c115 4 Vss 0.190935f
c116 2 Vss 0.189512f
r117 83 87 0.326018
r118 82 85 0.551426
r119 82 83 5.50157
r120 81 85 0.551426
r121 80 81 18.3386
r122 76 85 0.0828784
r123 76 78 1.82344
r124 74 80 0.652036
r125 74 75 10.1279
r126 72 98 1.16709
r127 70 75 0.652036
r128 70 72 2.16729
r129 69 84 0.494161
r130 68 87 0.326018
r131 68 69 13.0037
r132 64 84 0.128424
r133 64 66 6.16843
r134 62 84 0.494161
r135 62 63 7.46046
r136 60 89 1.16709
r137 58 63 0.652036
r138 58 60 2.16729
r139 56 78 1.16709
r140 52 66 1.16709
r141 44 98 0.0476429
r142 44 46 1.92555
r143 39 46 0.5835
r144 38 40 0.652036
r145 38 39 2.8008
r146 35 46 0.0685365
r147 31 89 0.0476429
r148 29 31 1.45875
r149 28 32 0.652036
r150 28 31 1.45875
r151 25 29 0.652036
r152 14 56 0.123773
r153 12 40 5.1348
r154 10 52 0.123773
r155 8 35 5.1348
r156 6 52 0.123773
r157 4 25 5.1348
r158 2 32 5.1348
.ends

.subckt PM_G3_MUXI2_N3_SELI 2 4 6 8 21 29 33 35 38 43 53 58 72 77 78 Vss
c62 78 Vss 8.12386e-19
c63 72 Vss 0.00203892f
c64 58 Vss 0.00238787f
c65 53 Vss 0.00260984f
c66 43 Vss 7.43568e-19
c67 38 Vss 0.00160083f
c68 36 Vss 0.00170119f
c69 35 Vss 0.00410624f
c70 33 Vss 0.00348196f
c71 29 Vss 0.00498872f
c72 21 Vss 0.166608f
c73 6 Vss 0.166608f
c74 4 Vss 0.00143493f
r75 77 78 0.655813
r76 76 77 3.501
r77 72 76 0.655813
r78 43 53 1.16709
r79 43 72 2.00578
r80 43 46 0.333429
r81 38 58 1.16709
r82 38 78 2.00578
r83 35 46 0.0685365
r84 35 36 7.46046
r85 31 36 0.652036
r86 31 33 7.91893
r87 29 33 1.16709
r88 21 58 0.50025
r89 18 53 0.50025
r90 8 21 4.37625
r91 6 18 4.37625
r92 4 29 0.123773
r93 2 29 0.123773
.ends

.subckt PM_G3_MUXI2_N3_SEL 2 4 6 8 16 22 26 37 40 42 46 51 58 63 68 72 77 78 Vss
c61 78 Vss 6.45399e-20
c62 77 Vss 9.69437e-20
c63 72 Vss 9.15408e-19
c64 68 Vss 0.00231917f
c65 63 Vss 0.00272254f
c66 58 Vss 0.00263414f
c67 51 Vss 5.38256e-19
c68 46 Vss 2.72603e-19
c69 42 Vss 0.00115861f
c70 37 Vss 0.00194091f
c71 26 Vss 0.166758f
c72 22 Vss 0.180313f
c73 20 Vss 0.0247918f
c74 17 Vss 0.0369697f
c75 16 Vss 0.191525f
c76 8 Vss 0.166608f
c77 2 Vss 0.193774f
r78 76 78 0.655813
r79 76 77 3.501
r80 72 77 0.655813
r81 54 63 1.16709
r82 54 72 2.00578
r83 51 54 0.5835
r84 49 58 1.16709
r85 46 49 0.5835
r86 42 68 1.16709
r87 42 78 2.00578
r88 38 46 0.0685365
r89 38 40 1.45875
r90 37 51 0.0685365
r91 37 40 3.12589
r92 36 58 0.0476429
r93 33 68 0.50025
r94 26 63 0.50025
r95 22 58 0.357321
r96 20 36 0.326018
r97 20 22 0.40845
r98 17 36 6.7686
r99 16 36 0.326018
r100 16 36 0.1167
r101 13 17 0.652036
r102 8 33 4.37625
r103 6 26 4.37625
r104 4 22 4.72635
r105 2 13 5.1348
.ends

.subckt PM_G3_MUXI2_N3_B 2 4 7 16 20 25 28 Vss
c23 28 Vss 0.00703355f
c24 25 Vss 5.28389e-19
c25 20 Vss 0.0287936f
c26 16 Vss 0.0658163f
c27 7 Vss 0.142278f
c28 4 Vss 0.40422f
c29 2 Vss 0.170892f
r30 22 28 1.16709
r31 22 25 0.0364688
r32 16 28 0.50025
r33 16 18 1.9839
r34 12 20 0.494161
r35 9 20 0.494161
r36 8 18 0.0685365
r37 7 20 0.128424
r38 7 8 4.7847
r39 4 12 12.3118
r40 2 9 4.49295
.ends

.subckt PM_G3_MUXI2_N3_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00389294f
c33 27 Vss 0.0072311f
c34 23 Vss 0.0072311f
c35 8 Vss 0.00143493f
c36 6 Vss 0.00143493f
r37 33 35 5.91836
r38 30 33 6.91864
r39 27 35 1.16709
r40 23 30 1.16709
r41 8 27 0.123773
r42 6 23 0.123773
r43 4 27 0.123773
r44 2 23 0.123773
.ends

.subckt PM_G3_MUXI2_N3_A 2 4 12 14 17 23 Vss
c24 23 Vss 0.00593108f
c25 17 Vss 2.08619e-19
c26 14 Vss 0.0835366f
c27 2 Vss 0.666088f
r28 20 23 1.16709
r29 17 20 0.0416786
r30 12 23 0.0476429
r31 12 14 1.92555
r32 7 14 0.0685365
r33 2 4 17.9718
r34 2 7 5.1348
.ends

.subckt G3_MUXI2_N3  VSS VDD SEL B Z A
*
* A	A
* Z	Z
* B	B
* SEL	SEL
* VDD	VDD
* VSS	VSS
XI12.X0 N_SELI_XI12.X0_D N_VDD_XI12.X0_PGD N_SEL_XI12.X0_CG N_VDD_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW12
XI13.X0 N_SELI_XI13.X0_D N_VSS_XI13.X0_PGD N_SEL_XI13.X0_CG N_VSS_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW12
XI17.X0 N_Z_XI17.X0_D N_VDD_XI17.X0_PGD N_SELI_XI17.X0_CG N_B_XI17.X0_PGS
+ N_VSS_XI17.X0_S TIGFET_HPNW12
XI15.X0 N_Z_XI15.X0_D N_VSS_XI15.X0_PGD N_SEL_XI15.X0_CG N_B_XI15.X0_PGS
+ N_VDD_XI15.X0_S TIGFET_HPNW12
XI16.X0 N_Z_XI16.X0_D N_VDD_XI16.X0_PGD N_SEL_XI16.X0_CG N_A_XI16.X0_PGS
+ N_VSS_XI16.X0_S TIGFET_HPNW12
XI14.X0 N_Z_XI14.X0_D N_VSS_XI14.X0_PGD N_SELI_XI14.X0_CG N_A_XI14.X0_PGS
+ N_VDD_XI14.X0_S TIGFET_HPNW12
*
x_PM_G3_MUXI2_N3_VSS N_VSS_XI12.X0_S N_VSS_XI13.X0_PGD N_VSS_XI13.X0_PGS
+ N_VSS_XI17.X0_S N_VSS_XI15.X0_PGD N_VSS_XI16.X0_S N_VSS_XI14.X0_PGD
+ N_VSS_c_4_p N_VSS_c_20_p N_VSS_c_44_p N_VSS_c_67_p N_VSS_c_69_p N_VSS_c_45_p
+ N_VSS_c_5_p N_VSS_c_26_p N_VSS_c_17_p N_VSS_c_27_p N_VSS_c_9_p N_VSS_c_19_p
+ N_VSS_c_6_p N_VSS_c_10_p N_VSS_c_11_p N_VSS_c_28_p N_VSS_c_24_p N_VSS_c_30_p
+ N_VSS_c_32_p N_VSS_c_33_p VSS N_VSS_c_12_p N_VSS_c_25_p N_VSS_c_34_p Vss
+ PM_G3_MUXI2_N3_VSS
x_PM_G3_MUXI2_N3_VDD N_VDD_XI12.X0_PGD N_VDD_XI12.X0_PGS N_VDD_XI13.X0_S
+ N_VDD_XI17.X0_PGD N_VDD_XI15.X0_S N_VDD_XI16.X0_PGD N_VDD_XI14.X0_S
+ N_VDD_c_81_n N_VDD_c_164_p N_VDD_c_128_p N_VDD_c_121_p N_VDD_c_144_p
+ N_VDD_c_82_n N_VDD_c_84_n N_VDD_c_90_n N_VDD_c_91_n N_VDD_c_97_n N_VDD_c_103_n
+ N_VDD_c_104_n N_VDD_c_106_n N_VDD_c_107_n N_VDD_c_108_n N_VDD_c_112_n
+ N_VDD_c_116_n N_VDD_c_117_n VDD N_VDD_c_118_n N_VDD_c_120_n Vss
+ PM_G3_MUXI2_N3_VDD
x_PM_G3_MUXI2_N3_SELI N_SELI_XI12.X0_D N_SELI_XI13.X0_D N_SELI_XI17.X0_CG
+ N_SELI_XI14.X0_CG N_SELI_c_229_p N_SELI_c_169_n N_SELI_c_171_n N_SELI_c_174_n
+ N_SELI_c_175_n N_SELI_c_188_n N_SELI_c_191_n N_SELI_c_178_n N_SELI_c_179_n
+ N_SELI_c_180_n N_SELI_c_211_p Vss PM_G3_MUXI2_N3_SELI
x_PM_G3_MUXI2_N3_SEL N_SEL_XI12.X0_CG N_SEL_XI13.X0_CG N_SEL_XI15.X0_CG
+ N_SEL_XI16.X0_CG N_SEL_c_231_n N_SEL_c_272_p N_SEL_c_273_p N_SEL_c_232_n SEL
+ N_SEL_c_233_n N_SEL_c_234_n N_SEL_c_257_n N_SEL_c_236_n N_SEL_c_260_n
+ N_SEL_c_246_n N_SEL_c_237_n N_SEL_c_239_n N_SEL_c_240_n Vss PM_G3_MUXI2_N3_SEL
x_PM_G3_MUXI2_N3_B N_B_XI17.X0_PGS N_B_XI15.X0_PGS N_B_c_292_n N_B_c_310_n
+ N_B_c_301_n B N_B_c_293_n Vss PM_G3_MUXI2_N3_B
x_PM_G3_MUXI2_N3_Z N_Z_XI17.X0_D N_Z_XI15.X0_D N_Z_XI16.X0_D N_Z_XI14.X0_D
+ N_Z_c_315_n N_Z_c_325_n N_Z_c_319_n Z Vss PM_G3_MUXI2_N3_Z
x_PM_G3_MUXI2_N3_A N_A_XI16.X0_PGS N_A_XI14.X0_PGS N_A_c_366_n N_A_c_350_n A
+ N_A_c_356_n Vss PM_G3_MUXI2_N3_A
cc_1 N_VSS_XI13.X0_PGD N_VDD_XI12.X0_PGD 0.00200584f
cc_2 N_VSS_XI15.X0_PGD N_VDD_XI17.X0_PGD 2.44446e-19
cc_3 N_VSS_XI14.X0_PGD N_VDD_XI16.X0_PGD 2.44446e-19
cc_4 N_VSS_c_4_p N_VDD_c_81_n 0.00200584f
cc_5 N_VSS_c_5_p N_VDD_c_82_n 9.64791e-19
cc_6 N_VSS_c_6_p N_VDD_c_82_n 4.10707e-19
cc_7 N_VSS_c_4_p N_VDD_c_84_n 3.89167e-19
cc_8 N_VSS_c_5_p N_VDD_c_84_n 0.00161703f
cc_9 N_VSS_c_9_p N_VDD_c_84_n 2.26455e-19
cc_10 N_VSS_c_10_p N_VDD_c_84_n 0.00442837f
cc_11 N_VSS_c_11_p N_VDD_c_84_n 0.00129625f
cc_12 N_VSS_c_12_p N_VDD_c_84_n 7.74609e-19
cc_13 N_VSS_c_10_p N_VDD_c_90_n 0.00157719f
cc_14 N_VSS_XI13.X0_PGS N_VDD_c_91_n 2.59535e-19
cc_15 N_VSS_XI15.X0_PGD N_VDD_c_91_n 2.19376e-19
cc_16 N_VSS_c_5_p N_VDD_c_91_n 0.00180638f
cc_17 N_VSS_c_17_p N_VDD_c_91_n 7.4365e-19
cc_18 N_VSS_c_9_p N_VDD_c_91_n 9.55109e-19
cc_19 N_VSS_c_19_p N_VDD_c_91_n 2.70301e-19
cc_20 N_VSS_c_20_p N_VDD_c_97_n 0.0011044f
cc_21 N_VSS_c_17_p N_VDD_c_97_n 0.00161703f
cc_22 N_VSS_c_19_p N_VDD_c_97_n 2.26455e-19
cc_23 N_VSS_c_11_p N_VDD_c_97_n 0.00590664f
cc_24 N_VSS_c_24_p N_VDD_c_97_n 0.0034989f
cc_25 N_VSS_c_25_p N_VDD_c_97_n 7.61747e-19
cc_26 N_VSS_c_26_p N_VDD_c_103_n 0.00121523f
cc_27 N_VSS_c_27_p N_VDD_c_104_n 3.5277e-19
cc_28 N_VSS_c_28_p N_VDD_c_104_n 0.00873112f
cc_29 N_VSS_c_28_p N_VDD_c_106_n 0.00155968f
cc_30 N_VSS_c_30_p N_VDD_c_107_n 4.01154e-19
cc_31 N_VSS_c_27_p N_VDD_c_108_n 0.00187494f
cc_32 N_VSS_c_32_p N_VDD_c_108_n 0.0041789f
cc_33 N_VSS_c_33_p N_VDD_c_108_n 0.0078367f
cc_34 N_VSS_c_34_p N_VDD_c_108_n 9.16632e-19
cc_35 N_VSS_c_17_p N_VDD_c_112_n 4.28751e-19
cc_36 N_VSS_c_19_p N_VDD_c_112_n 6.0691e-19
cc_37 N_VSS_c_24_p N_VDD_c_112_n 0.00108024f
cc_38 N_VSS_c_33_p N_VDD_c_112_n 0.00418449f
cc_39 N_VSS_c_11_p N_VDD_c_116_n 0.00121059f
cc_40 N_VSS_c_33_p N_VDD_c_117_n 0.00100712f
cc_41 N_VSS_c_5_p N_VDD_c_118_n 3.48267e-19
cc_42 N_VSS_c_9_p N_VDD_c_118_n 6.46219e-19
cc_43 N_VSS_c_26_p N_VDD_c_120_n 2.82095e-19
cc_44 N_VSS_c_44_p N_SELI_c_169_n 3.43419e-19
cc_45 N_VSS_c_45_p N_SELI_c_169_n 3.48267e-19
cc_46 N_VSS_c_44_p N_SELI_c_171_n 3.48267e-19
cc_47 N_VSS_c_45_p N_SELI_c_171_n 8.50248e-19
cc_48 N_VSS_c_10_p N_SELI_c_171_n 2.24858e-19
cc_49 N_VSS_c_26_p N_SELI_c_174_n 7.64616e-19
cc_50 N_VSS_c_17_p N_SELI_c_175_n 2.2375e-19
cc_51 N_VSS_c_19_p N_SELI_c_175_n 2.18171e-19
cc_52 N_VSS_c_33_p N_SELI_c_175_n 9.07743e-19
cc_53 N_VSS_c_17_p N_SELI_c_178_n 2.15082e-19
cc_54 N_VSS_c_28_p N_SELI_c_179_n 5.93394e-19
cc_55 N_VSS_c_33_p N_SELI_c_180_n 5.03655e-19
cc_56 N_VSS_XI13.X0_PGD N_SEL_c_231_n 4.23684e-19
cc_57 N_VSS_c_11_p N_SEL_c_232_n 4.38015e-19
cc_58 N_VSS_c_33_p N_SEL_c_233_n 7.91494e-19
cc_59 N_VSS_c_5_p N_SEL_c_234_n 2.10271e-19
cc_60 N_VSS_c_9_p N_SEL_c_234_n 2.26251e-19
cc_61 N_VSS_c_5_p N_SEL_c_236_n 2.15082e-19
cc_62 N_VSS_c_11_p N_SEL_c_237_n 7.83225e-19
cc_63 N_VSS_c_28_p N_SEL_c_237_n 2.12674e-19
cc_64 N_VSS_c_33_p N_SEL_c_239_n 4.36463e-19
cc_65 N_VSS_c_28_p N_SEL_c_240_n 7.26277e-19
cc_66 N_VSS_XI13.X0_PGS N_B_c_292_n 2.57132e-19
cc_67 N_VSS_c_67_p N_B_c_293_n 0.00132057f
cc_68 N_VSS_c_67_p N_Z_c_315_n 3.43419e-19
cc_69 N_VSS_c_69_p N_Z_c_315_n 3.43419e-19
cc_70 N_VSS_c_26_p N_Z_c_315_n 3.48267e-19
cc_71 N_VSS_c_27_p N_Z_c_315_n 3.48267e-19
cc_72 N_VSS_c_67_p N_Z_c_319_n 3.48267e-19
cc_73 N_VSS_c_69_p N_Z_c_319_n 3.48267e-19
cc_74 N_VSS_c_26_p N_Z_c_319_n 5.68482e-19
cc_75 N_VSS_c_27_p N_Z_c_319_n 5.71987e-19
cc_76 N_VSS_c_33_p N_Z_c_319_n 9.78034e-19
cc_77 N_VSS_c_28_p A 2.12185e-19
cc_78 N_VDD_c_121_p N_SELI_c_169_n 3.43419e-19
cc_79 N_VDD_c_84_n N_SELI_c_169_n 2.74986e-19
cc_80 N_VDD_c_91_n N_SELI_c_169_n 3.48267e-19
cc_81 N_VDD_c_121_p N_SELI_c_171_n 3.48267e-19
cc_82 N_VDD_c_84_n N_SELI_c_171_n 3.83029e-19
cc_83 N_VDD_c_91_n N_SELI_c_171_n 7.09569e-19
cc_84 N_VDD_c_108_n N_SELI_c_175_n 6.15494e-19
cc_85 N_VDD_c_128_p N_SELI_c_188_n 2.21762e-19
cc_86 N_VDD_c_103_n N_SELI_c_188_n 2.87975e-19
cc_87 N_VDD_c_120_n N_SELI_c_188_n 2.30774e-19
cc_88 N_VDD_c_103_n N_SELI_c_191_n 2.28697e-19
cc_89 N_VDD_c_108_n N_SELI_c_178_n 3.66936e-19
cc_90 N_VDD_XI12.X0_PGD N_SEL_c_231_n 4.31283e-19
cc_91 N_VDD_c_121_p N_SEL_c_232_n 4.75243e-19
cc_92 N_VDD_c_91_n N_SEL_c_232_n 8.22147e-19
cc_93 N_VDD_c_104_n N_SEL_c_233_n 2.47222e-19
cc_94 N_VDD_c_108_n N_SEL_c_233_n 6.15494e-19
cc_95 N_VDD_c_108_n N_SEL_c_246_n 3.66936e-19
cc_96 N_VDD_c_97_n N_SEL_c_237_n 3.65289e-19
cc_97 N_VDD_c_108_n N_SEL_c_239_n 2.2501e-19
cc_98 N_VDD_c_121_p N_B_c_292_n 2.35559e-19
cc_99 N_VDD_c_104_n N_Z_c_315_n 2.74986e-19
cc_100 N_VDD_c_121_p N_Z_c_325_n 3.43419e-19
cc_101 N_VDD_c_144_p N_Z_c_325_n 3.43419e-19
cc_102 N_VDD_c_91_n N_Z_c_325_n 3.48267e-19
cc_103 N_VDD_c_97_n N_Z_c_325_n 2.74986e-19
cc_104 N_VDD_c_107_n N_Z_c_325_n 3.72199e-19
cc_105 N_VDD_c_121_p N_Z_c_319_n 3.48267e-19
cc_106 N_VDD_c_144_p N_Z_c_319_n 3.48267e-19
cc_107 N_VDD_c_91_n N_Z_c_319_n 8.16241e-19
cc_108 N_VDD_c_97_n N_Z_c_319_n 3.83904e-19
cc_109 N_VDD_c_104_n N_Z_c_319_n 3.83904e-19
cc_110 N_VDD_c_107_n N_Z_c_319_n 8.08807e-19
cc_111 N_VDD_c_108_n N_Z_c_319_n 0.00135474f
cc_112 N_VDD_XI16.X0_PGD N_A_XI16.X0_PGS 0.00146246f
cc_113 N_VDD_c_108_n N_A_XI16.X0_PGS 0.00109285f
cc_114 N_VDD_c_104_n N_A_c_350_n 3.5103e-19
cc_115 N_VDD_c_108_n N_A_c_350_n 3.92527e-19
cc_116 N_VDD_c_103_n A 5.27373e-19
cc_117 N_VDD_c_104_n A 0.00141439f
cc_118 N_VDD_c_108_n A 5.06354e-19
cc_119 N_VDD_c_120_n A 3.44698e-19
cc_120 N_VDD_XI16.X0_PGD N_A_c_356_n 3.32271e-19
cc_121 N_VDD_c_164_p N_A_c_356_n 0.00480616f
cc_122 N_VDD_c_103_n N_A_c_356_n 3.95721e-19
cc_123 N_VDD_c_104_n N_A_c_356_n 0.00120343f
cc_124 N_VDD_c_108_n N_A_c_356_n 3.70842e-19
cc_125 N_VDD_c_120_n N_A_c_356_n 6.02643e-19
cc_126 N_SELI_c_169_n N_SEL_c_231_n 7.69306e-19
cc_127 N_SELI_c_171_n N_SEL_c_231_n 9.27181e-19
cc_128 N_SELI_c_174_n N_SEL_c_231_n 4.0622e-19
cc_129 N_SELI_c_188_n N_SEL_c_232_n 0.00290285f
cc_130 N_SELI_c_175_n N_SEL_c_233_n 0.00242961f
cc_131 N_SELI_c_178_n N_SEL_c_233_n 4.99367e-19
cc_132 N_SELI_c_171_n N_SEL_c_234_n 0.0024269f
cc_133 N_SELI_c_174_n N_SEL_c_234_n 0.00290285f
cc_134 N_SELI_c_191_n N_SEL_c_257_n 5.42085e-19
cc_135 N_SELI_c_171_n N_SEL_c_236_n 0.00100994f
cc_136 N_SELI_c_174_n N_SEL_c_236_n 5.63096e-19
cc_137 N_SELI_c_191_n N_SEL_c_260_n 0.00494389f
cc_138 N_SELI_c_178_n N_SEL_c_260_n 8.7809e-19
cc_139 N_SELI_c_191_n N_SEL_c_246_n 8.69867e-19
cc_140 N_SELI_c_178_n N_SEL_c_246_n 0.00494884f
cc_141 N_SELI_c_175_n N_SEL_c_237_n 0.00165721f
cc_142 N_SELI_c_188_n N_SEL_c_237_n 4.7869e-19
cc_143 N_SELI_c_179_n N_SEL_c_237_n 9.92651e-19
cc_144 N_SELI_c_211_p N_SEL_c_237_n 8.15293e-19
cc_145 N_SELI_c_171_n N_SEL_c_239_n 3.01017e-19
cc_146 N_SELI_c_180_n N_SEL_c_239_n 0.00144491f
cc_147 N_SELI_c_188_n N_SEL_c_240_n 0.00165436f
cc_148 N_SELI_c_179_n N_SEL_c_240_n 8.14736e-19
cc_149 N_SELI_XI17.X0_CG N_B_XI17.X0_PGS 4.31731e-19
cc_150 N_SELI_c_191_n N_B_XI17.X0_PGS 6.66106e-19
cc_151 N_SELI_c_171_n N_B_XI15.X0_PGS 2.97793e-19
cc_152 N_SELI_c_174_n N_B_XI15.X0_PGS 3.99745e-19
cc_153 N_SELI_c_191_n N_B_XI15.X0_PGS 5.45575e-19
cc_154 N_SELI_c_174_n N_B_c_292_n 4.07501e-19
cc_155 N_SELI_c_174_n N_B_c_301_n 5.40503e-19
cc_156 N_SELI_c_191_n N_B_c_301_n 0.00179467f
cc_157 N_SELI_c_174_n B 0.0012894f
cc_158 N_SELI_c_174_n N_B_c_293_n 0.00106912f
cc_159 N_SELI_c_171_n N_Z_c_319_n 0.00105053f
cc_160 N_SELI_c_175_n N_Z_c_319_n 0.00208341f
cc_161 N_SELI_c_188_n N_Z_c_319_n 0.00213869f
cc_162 N_SELI_c_229_p N_A_XI16.X0_PGS 4.87172e-19
cc_163 N_SELI_c_178_n N_A_XI16.X0_PGS 0.00276355f
cc_164 N_SEL_c_272_p N_B_XI15.X0_PGS 2.04953e-19
cc_165 N_SEL_c_273_p N_B_XI15.X0_PGS 4.65537e-19
cc_166 N_SEL_c_232_n N_B_XI15.X0_PGS 8.40923e-19
cc_167 N_SEL_c_236_n N_B_XI15.X0_PGS 0.00100354f
cc_168 N_SEL_c_260_n N_B_XI15.X0_PGS 0.00202689f
cc_169 N_SEL_c_232_n N_B_c_310_n 2.88938e-19
cc_170 N_SEL_c_236_n N_B_c_310_n 7.65159e-19
cc_171 N_SEL_c_236_n N_B_c_293_n 0.00115283f
cc_172 N_SEL_c_233_n N_Z_c_319_n 0.00189968f
cc_173 N_SEL_c_257_n N_Z_c_319_n 0.00240311f
cc_174 N_SEL_c_246_n N_Z_c_319_n 9.35582e-19
cc_175 N_SEL_c_237_n N_Z_c_319_n 9.65156e-19
cc_176 N_SEL_c_239_n N_Z_c_319_n 0.0021646f
cc_177 N_SEL_c_240_n N_Z_c_319_n 9.51045e-19
cc_178 N_SEL_XI16.X0_CG N_A_XI16.X0_PGS 4.87172e-19
cc_179 N_SEL_c_246_n N_A_XI16.X0_PGS 0.00276355f
cc_180 N_SEL_c_233_n N_A_c_366_n 2.18171e-19
cc_181 N_SEL_c_233_n A 2.78876e-19
cc_182 N_SEL_c_246_n A 2.15082e-19
cc_183 N_SEL_c_233_n N_A_c_356_n 2.30774e-19
cc_184 B N_Z_c_319_n 4.05731e-19
cc_185 N_B_XI17.X0_PGS N_A_XI16.X0_PGS 0.00134199f
*
.ends
*
*
.subckt MUXI2_HPNW12 A B S0 Y VDD VSS
xgate (VSS VDD S0 B Y A) G3_MUXI2_N3
.ends
*
* File: G2_NAND2_N3.pex.netlist
* Created: Sun Apr 10 19:03:25 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NAND2_N3_VSS 2 4 6 8 10 20 21 41 45 50 59 66 71 72 Vss
c25 72 Vss 8.04097e-19
c26 71 Vss 0.00222754f
c27 67 Vss 0.00133588f
c28 66 Vss 0.0113624f
c29 59 Vss 0.0053595f
c30 50 Vss 0.00153395f
c31 45 Vss 0.00130895f
c32 41 Vss 0.00965443f
c33 38 Vss 0.0299311f
c34 37 Vss 0.0299311f
c35 32 Vss 0.106916f
c36 27 Vss 0.0688416f
c37 21 Vss 0.0350852f
c38 20 Vss 0.0646396f
c39 10 Vss 0.190769f
c40 8 Vss 0.19123f
c41 6 Vss 0.189919f
c42 4 Vss 0.191018f
r43 71 73 0.652036
r44 71 72 4.33457
r45 64 72 0.652036
r46 64 66 12.5452
r47 63 67 0.655813
r48 63 66 6.50186
r49 50 59 1.16709
r50 50 73 2.16729
r51 45 67 1.82344
r52 41 45 1.16709
r53 33 38 0.494161
r54 32 34 0.652036
r55 32 33 2.9175
r56 29 38 0.128424
r57 28 37 0.494161
r58 27 38 0.494161
r59 27 28 2.8008
r60 24 37 0.128424
r61 23 59 0.0476429
r62 21 23 1.4004
r63 20 37 0.494161
r64 20 23 1.5171
r65 17 21 0.652036
r66 10 34 5.1348
r67 8 29 5.1348
r68 6 17 5.1348
r69 4 24 5.1348
r70 2 41 0.123773
.ends

.subckt PM_G2_NAND2_N3_VDD 2 4 6 15 17 22 27 30 31 33 35 36 37 41 46 48 51 57
+ Vss
c42 57 Vss 0.00431501f
c43 49 Vss 7.68513e-19
c44 48 Vss 0.00721617f
c45 46 Vss 0.00728738f
c46 41 Vss 0.00103469f
c47 37 Vss 0.0066476f
c48 36 Vss 8.606e-19
c49 35 Vss 0.0118736f
c50 33 Vss 0.00172072f
c51 31 Vss 7.81221e-19
c52 30 Vss 0.00275683f
c53 27 Vss 0.00946889f
c54 22 Vss 0.00810168f
c55 17 Vss 0.170588f
c56 15 Vss 0.0352333f
c57 2 Vss 0.220859f
r58 48 51 0.326018
r59 47 49 0.551426
r60 47 48 5.37654
r61 46 49 0.551426
r62 45 46 8.41907
r63 43 64 1.16709
r64 41 49 0.0828784
r65 41 43 1.53169
r66 39 57 1.16709
r67 37 45 0.655813
r68 37 39 4.0845
r69 35 51 0.326018
r70 35 36 15.3377
r71 31 33 1.82344
r72 30 36 0.652036
r73 29 31 0.655813
r74 29 30 5.50157
r75 27 64 0.15
r76 22 33 1.16709
r77 17 57 0.428786
r78 15 17 5.3682
r79 12 15 0.652036
r80 6 27 0.123773
r81 4 22 0.123773
r82 2 12 6.3018
.ends

.subckt PM_G2_NAND2_N3_A 1 2 20 23 28 33 Vss
c18 33 Vss 0.00403439f
c19 28 Vss 0.00239607f
c20 20 Vss 0.0017793f
c21 12 Vss 0.166936f
c22 1 Vss 0.171396f
r23 25 33 1.16709
r24 23 25 3.00086
r25 20 28 1.16709
r26 20 23 2.37568
r27 12 33 0.50025
r28 9 28 0.50025
r29 2 12 4.37625
r30 1 9 4.60965
.ends

.subckt PM_G2_NAND2_N3_Z 2 4 6 18 22 25 28 Vss
c26 25 Vss 0.00178689f
c27 22 Vss 0.0056591f
c28 18 Vss 0.00911019f
c29 6 Vss 0.00143493f
r30 30 39 1.16709
r31 28 30 6.54354
r32 25 28 7.12704
r33 22 39 0.15
r34 18 25 1.16709
r35 6 22 0.123773
r36 4 22 0.123773
r37 2 18 0.123773
.ends

.subckt PM_G2_NAND2_N3_B 2 3 9 10 13 19 Vss
c23 19 Vss 1.07412e-19
c24 13 Vss 0.244723f
c25 10 Vss 0.0357412f
c26 9 Vss 0.288308f
c27 2 Vss 0.328264f
r28 19 22 0.125036
r29 13 22 1.16709
r30 11 13 2.39235
r31 9 11 0.652036
r32 9 10 8.92755
r33 6 10 0.652036
r34 3 13 5.6016
r35 2 6 9.8028
.ends

.subckt G2_NAND2_N3  VSS VDD A Z B
*
* B	B
* Z	Z
* A	A
* VDD	VDD
* VSS	VSS
XI13.X0 N_Z_XI13.X0_D N_VDD_XI13.X0_PGD N_A_XI13.X0_CG N_B_XI13.X0_PGS
+ N_VSS_XI13.X0_S TIGFET_HPNW12
XI14.X0 N_Z_XI14.X0_D N_VSS_XI14.X0_PGD N_A_XI14.X0_CG N_VSS_XI14.X0_PGS
+ N_VDD_XI14.X0_S TIGFET_HPNW12
XI15.X0 N_Z_XI15.X0_D N_VSS_XI15.X0_PGD N_B_XI15.X0_CG N_VSS_XI15.X0_PGS
+ N_VDD_XI15.X0_S TIGFET_HPNW12
*
x_PM_G2_NAND2_N3_VSS N_VSS_XI13.X0_S N_VSS_XI14.X0_PGD N_VSS_XI14.X0_PGS
+ N_VSS_XI15.X0_PGD N_VSS_XI15.X0_PGS N_VSS_c_6_p N_VSS_c_7_p N_VSS_c_19_p
+ N_VSS_c_5_p N_VSS_c_2_p N_VSS_c_9_p VSS N_VSS_c_10_p N_VSS_c_11_p Vss
+ PM_G2_NAND2_N3_VSS
x_PM_G2_NAND2_N3_VDD N_VDD_XI13.X0_PGD N_VDD_XI14.X0_S N_VDD_XI15.X0_S
+ N_VDD_c_60_p N_VDD_c_50_p N_VDD_c_44_p N_VDD_c_45_p N_VDD_c_26_n N_VDD_c_29_n
+ N_VDD_c_30_n N_VDD_c_31_n N_VDD_c_36_n N_VDD_c_55_p N_VDD_c_48_p N_VDD_c_41_p
+ N_VDD_c_37_n VDD N_VDD_c_43_p Vss PM_G2_NAND2_N3_VDD
x_PM_G2_NAND2_N3_A N_A_XI13.X0_CG N_A_XI14.X0_CG N_A_c_68_n A N_A_c_74_n
+ N_A_c_70_n Vss PM_G2_NAND2_N3_A
x_PM_G2_NAND2_N3_Z N_Z_XI13.X0_D N_Z_XI14.X0_D N_Z_XI15.X0_D N_Z_c_86_n
+ N_Z_c_90_n N_Z_c_88_n Z Vss PM_G2_NAND2_N3_Z
x_PM_G2_NAND2_N3_B N_B_XI13.X0_PGS N_B_XI15.X0_CG N_B_c_112_n N_B_c_114_n
+ N_B_c_117_n B Vss PM_G2_NAND2_N3_B
cc_1 N_VSS_XI14.X0_PGS N_VDD_c_26_n 3.44373e-19
cc_2 N_VSS_c_2_p N_VDD_c_26_n 4.83895e-19
cc_3 VSS N_VDD_c_26_n 0.00361022f
cc_4 VSS N_VDD_c_29_n 0.00159527f
cc_5 N_VSS_c_5_p N_VDD_c_30_n 3.7872e-19
cc_6 N_VSS_c_6_p N_VDD_c_31_n 0.00194111f
cc_7 N_VSS_c_7_p N_VDD_c_31_n 3.76573e-19
cc_8 N_VSS_c_2_p N_VDD_c_31_n 0.00161703f
cc_9 N_VSS_c_9_p N_VDD_c_31_n 2.26455e-19
cc_10 N_VSS_c_10_p N_VDD_c_31_n 0.00519315f
cc_11 N_VSS_c_11_p N_VDD_c_36_n 0.00104854f
cc_12 N_VSS_XI15.X0_PGS N_VDD_c_37_n 4.24059e-19
cc_13 N_VSS_c_2_p N_VDD_c_37_n 5.47905e-19
cc_14 VSS N_VDD_c_37_n 2.38209e-19
cc_15 N_VSS_c_9_p N_A_c_68_n 2.354e-19
cc_16 VSS N_A_c_68_n 0.00258255f
cc_17 N_VSS_c_2_p N_A_c_70_n 2.15082e-19
cc_18 N_VSS_c_9_p N_A_c_70_n 4.9359e-19
cc_19 N_VSS_c_19_p N_Z_c_86_n 3.43419e-19
cc_20 N_VSS_c_5_p N_Z_c_86_n 3.48267e-19
cc_21 N_VSS_c_5_p N_Z_c_88_n 8.92744e-19
cc_22 VSS N_Z_c_88_n 0.0013442f
cc_23 N_VSS_XI14.X0_PGD N_B_c_112_n 7.63854e-19
cc_24 N_VSS_XI15.X0_PGD N_B_c_112_n 7.63854e-19
cc_25 N_VSS_XI14.X0_PGS N_B_c_114_n 9.45978e-19
cc_26 N_VDD_XI13.X0_PGD N_A_XI13.X0_CG 4.9269e-19
cc_27 N_VDD_c_41_p N_A_c_68_n 2.11067e-19
cc_28 N_VDD_XI13.X0_PGD N_A_c_74_n 4.86892e-19
cc_29 N_VDD_c_43_p N_A_c_74_n 5.00305e-19
cc_30 N_VDD_c_44_p N_Z_c_90_n 3.43419e-19
cc_31 N_VDD_c_45_p N_Z_c_90_n 3.43419e-19
cc_32 N_VDD_c_30_n N_Z_c_90_n 3.72199e-19
cc_33 N_VDD_c_31_n N_Z_c_90_n 2.82909e-19
cc_34 N_VDD_c_48_p N_Z_c_90_n 3.70313e-19
cc_35 N_VDD_XI13.X0_PGD N_Z_c_88_n 3.98301e-19
cc_36 N_VDD_c_50_p N_Z_c_88_n 6.23961e-19
cc_37 N_VDD_c_44_p N_Z_c_88_n 3.48267e-19
cc_38 N_VDD_c_45_p N_Z_c_88_n 3.48267e-19
cc_39 N_VDD_c_30_n N_Z_c_88_n 8.08807e-19
cc_40 N_VDD_c_31_n N_Z_c_88_n 5.69519e-19
cc_41 N_VDD_c_55_p N_Z_c_88_n 0.00170631f
cc_42 N_VDD_c_48_p N_Z_c_88_n 8.48488e-19
cc_43 N_VDD_c_41_p N_Z_c_88_n 0.00275333f
cc_44 N_VDD_c_43_p N_Z_c_88_n 9.31683e-19
cc_45 N_VDD_XI13.X0_PGD N_B_XI13.X0_PGS 0.00331576f
cc_46 N_VDD_c_60_p N_B_c_112_n 0.00812117f
cc_47 N_VDD_c_55_p N_B_c_117_n 3.69683e-19
cc_48 N_VDD_c_41_p N_B_c_117_n 6.28222e-19
cc_49 N_VDD_c_43_p N_B_c_117_n 0.00146481f
cc_50 N_VDD_c_31_n B 2.63427e-19
cc_51 N_VDD_c_55_p B 5.03854e-19
cc_52 N_VDD_c_41_p B 7.0924e-19
cc_53 N_VDD_c_43_p B 3.69683e-19
cc_54 N_A_c_68_n N_Z_c_88_n 0.00825864f
cc_55 N_A_c_74_n N_Z_c_88_n 8.85473e-19
cc_56 N_A_c_70_n N_Z_c_88_n 0.00100714f
cc_57 N_A_XI13.X0_CG N_B_XI13.X0_PGS 4.97429e-19
cc_58 N_A_c_68_n N_B_XI13.X0_PGS 5.60962e-19
cc_59 N_A_c_74_n N_B_XI13.X0_PGS 5.64689e-19
cc_60 N_A_c_68_n N_B_c_112_n 3.152e-19
cc_61 N_A_c_74_n N_B_c_112_n 7.5465e-19
cc_62 N_A_c_70_n N_B_c_112_n 0.00132909f
cc_63 N_A_c_70_n N_B_c_117_n 9.27569e-19
cc_64 N_Z_c_90_n N_B_c_112_n 3.31584e-19
cc_65 N_Z_c_88_n N_B_c_112_n 4.20335e-19
cc_66 N_Z_c_88_n N_B_c_117_n 0.00101313f
cc_67 N_Z_c_88_n B 0.00147455f
*
.ends
*
*
.subckt NAND2_HPNW12 A B Y VDD VSS
xgate (VSS VDD A Y B) G2_NAND2_N3
.ends
*
* File: G2_NOR2_N3.pex.netlist
* Created: Mon Feb 28 10:13:32 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NOR2_N3_VSS 2 4 6 18 23 28 31 36 41 50 59 60 64 65 70 73 74 79 Vss
c39 74 Vss 3.75522e-19
c40 73 Vss 0.0047697f
c41 70 Vss 0.00562567f
c42 65 Vss 8.27694e-19
c43 64 Vss 0.00178035f
c44 60 Vss 6.04131e-19
c45 59 Vss 0.00565031f
c46 50 Vss 0.00520705f
c47 41 Vss 0.00279442f
c48 36 Vss 0.00113197f
c49 31 Vss 0.00124387f
c50 28 Vss 0.00807325f
c51 23 Vss 0.00817292f
c52 18 Vss 0.089128f
c53 4 Vss 0.189873f
r54 73 79 0.326018
r55 72 77 0.14525
r56 72 73 5.50157
r57 71 74 0.494161
r58 70 79 0.326018
r59 70 71 10.1279
r60 66 74 0.128424
r61 64 74 0.494161
r62 64 65 4.37625
r63 59 65 0.652036
r64 58 60 0.655813
r65 58 59 18.3386
r66 41 77 2.334
r67 36 50 1.16709
r68 36 66 2.16729
r69 31 60 1.82344
r70 28 41 1.16709
r71 23 31 1.16709
r72 16 50 0.0476429
r73 16 18 2.04225
r74 12 18 0.0685365
r75 6 28 0.123773
r76 4 12 5.1348
r77 2 23 0.123773
.ends

.subckt PM_G2_NOR2_N3_VDD 2 4 6 8 10 27 36 41 45 47 48 52 54 55 58 60 62 64 66
+ 72 78 Vss
c45 78 Vss 0.00622884f
c46 72 Vss 0.00491473f
c47 64 Vss 4.52364e-19
c48 62 Vss 0.00102348f
c49 60 Vss 6.08701e-19
c50 58 Vss 0.00198853f
c51 55 Vss 8.64913e-19
c52 54 Vss 0.00550278f
c53 52 Vss 0.0017471f
c54 49 Vss 0.0017501f
c55 48 Vss 0.00518267f
c56 47 Vss 0.00321334f
c57 45 Vss 0.0127334f
c58 41 Vss 0.00818763f
c59 37 Vss 0.129193f
c60 36 Vss 7.7089e-20
c61 27 Vss 0.0356247f
c62 26 Vss 0.102427f
c63 10 Vss 0.190932f
c64 8 Vss 0.189362f
c65 4 Vss 0.190692f
c66 2 Vss 0.191746f
r67 72 75 0.05
r68 62 78 1.16709
r69 60 66 0.326018
r70 60 62 2.16729
r71 58 75 1.16709
r72 56 58 2.95918
r73 54 66 0.326018
r74 54 55 10.1696
r75 50 64 0.0828784
r76 50 52 1.82344
r77 48 56 0.652036
r78 48 49 4.37625
r79 47 55 0.652036
r80 46 64 0.551426
r81 46 47 5.50157
r82 45 64 0.551426
r83 44 49 0.652036
r84 44 45 19.0888
r85 41 52 1.16709
r86 36 72 0.0238214
r87 36 37 2.26917
r88 33 36 2.26917
r89 29 78 0.0476429
r90 27 29 1.5171
r91 26 30 0.652036
r92 26 29 1.4004
r93 23 27 0.652036
r94 20 37 0.00605528
r95 17 33 0.00605528
r96 10 30 5.1348
r97 8 23 5.1348
r98 6 41 0.123773
r99 4 17 5.1348
r100 2 20 5.1348
.ends

.subckt PM_G2_NOR2_N3_B 2 4 10 13 18 21 26 31 Vss
c20 31 Vss 0.0033745f
c21 26 Vss 0.00378619f
c22 18 Vss 0.00118409f
c23 13 Vss 0.166574f
c24 10 Vss 7.77222e-20
c25 2 Vss 0.16675f
r26 23 31 1.16709
r27 21 23 2.37568
r28 18 26 1.16709
r29 18 21 2.45904
r30 13 31 0.50025
r31 10 26 0.50025
r32 4 13 4.37625
r33 2 10 4.37625
.ends

.subckt PM_G2_NOR2_N3_Z 2 4 6 18 22 25 28 Vss
c24 25 Vss 0.00353787f
c25 22 Vss 0.0056593f
c26 18 Vss 0.00813452f
c27 6 Vss 0.00143493f
r28 28 30 6.16843
r29 25 28 6.66857
r30 22 30 1.16709
r31 18 25 1.16709
r32 6 22 0.123773
r33 4 22 0.123773
r34 2 18 0.123773
.ends

.subckt PM_G2_NOR2_N3_A 2 4 10 11 14 18 21 Vss
c18 18 Vss 2.27081e-19
c19 14 Vss 0.2392f
c20 11 Vss 0.0348811f
c21 10 Vss 0.282285f
c22 2 Vss 0.269802f
r23 18 27 1.16709
r24 18 21 0.0416786
r25 14 27 0.05
r26 12 14 2.27565
r27 10 12 0.652036
r28 10 11 8.92755
r29 7 11 0.652036
r30 4 14 5.6016
r31 2 7 7.87725
.ends

.subckt G2_NOR2_N3  VSS VDD B Z A
*
* A	A
* Z	Z
* B	B
* VDD	VDD
* VSS	VSS
XI8.X0 N_Z_XI8.X0_D N_VDD_XI8.X0_PGD N_B_XI8.X0_CG N_VDD_XI8.X0_PGS
+ N_VSS_XI8.X0_S TIGFET_HPNW12
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_A_XI6.X0_PGS N_VDD_XI6.X0_S
+ TIGFET_HPNW12
XI7.X0 N_Z_XI7.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW12
*
x_PM_G2_NOR2_N3_VSS N_VSS_XI8.X0_S N_VSS_XI6.X0_PGD N_VSS_XI7.X0_S N_VSS_c_2_p
+ N_VSS_c_8_p N_VSS_c_31_p N_VSS_c_3_p N_VSS_c_6_p N_VSS_c_32_p N_VSS_c_13_p
+ N_VSS_c_4_p N_VSS_c_5_p N_VSS_c_14_p N_VSS_c_17_p N_VSS_c_15_p N_VSS_c_20_p
+ N_VSS_c_16_p VSS Vss PM_G2_NOR2_N3_VSS
x_PM_G2_NOR2_N3_VDD N_VDD_XI8.X0_PGD N_VDD_XI8.X0_PGS N_VDD_XI6.X0_S
+ N_VDD_XI7.X0_PGD N_VDD_XI7.X0_PGS N_VDD_c_41_n N_VDD_c_63_p N_VDD_c_70_p
+ N_VDD_c_42_n N_VDD_c_45_n N_VDD_c_47_n N_VDD_c_49_n N_VDD_c_50_n N_VDD_c_56_n
+ N_VDD_c_65_p N_VDD_c_57_n N_VDD_c_58_n N_VDD_c_60_n VDD N_VDD_c_66_p
+ N_VDD_c_61_n Vss PM_G2_NOR2_N3_VDD
x_PM_G2_NOR2_N3_B N_B_XI8.X0_CG N_B_XI6.X0_CG N_B_c_90_n N_B_c_100_p N_B_c_85_n
+ B N_B_c_94_n N_B_c_88_n Vss PM_G2_NOR2_N3_B
x_PM_G2_NOR2_N3_Z N_Z_XI8.X0_D N_Z_XI6.X0_D N_Z_XI7.X0_D N_Z_c_105_n N_Z_c_107_n
+ N_Z_c_109_n Z Vss PM_G2_NOR2_N3_Z
x_PM_G2_NOR2_N3_A N_A_XI6.X0_PGS N_A_XI7.X0_CG N_A_c_129_n N_A_c_132_n
+ N_A_c_134_n N_A_c_136_n A Vss PM_G2_NOR2_N3_A
cc_1 N_VSS_XI6.X0_PGD N_VDD_XI7.X0_PGD 0.00209072f
cc_2 N_VSS_c_2_p N_VDD_c_41_n 0.00209072f
cc_3 N_VSS_c_3_p N_VDD_c_42_n 0.00187494f
cc_4 N_VSS_c_4_p N_VDD_c_42_n 0.00752502f
cc_5 N_VSS_c_5_p N_VDD_c_42_n 0.00189882f
cc_6 N_VSS_c_6_p N_VDD_c_45_n 4.76491e-19
cc_7 N_VSS_c_4_p N_VDD_c_45_n 0.00426824f
cc_8 N_VSS_c_8_p N_VDD_c_47_n 2.3316e-19
cc_9 N_VSS_c_3_p N_VDD_c_47_n 7.26139e-19
cc_10 N_VSS_c_3_p N_VDD_c_49_n 4.01154e-19
cc_11 N_VSS_c_2_p N_VDD_c_50_n 3.71132e-19
cc_12 N_VSS_c_6_p N_VDD_c_50_n 0.00141228f
cc_13 N_VSS_c_13_p N_VDD_c_50_n 0.00114511f
cc_14 N_VSS_c_14_p N_VDD_c_50_n 0.00352847f
cc_15 N_VSS_c_15_p N_VDD_c_50_n 0.00446295f
cc_16 N_VSS_c_16_p N_VDD_c_50_n 7.74609e-19
cc_17 N_VSS_c_17_p N_VDD_c_56_n 0.00106582f
cc_18 N_VSS_c_15_p N_VDD_c_57_n 0.00151536f
cc_19 N_VSS_c_6_p N_VDD_c_58_n 0.00109227f
cc_20 N_VSS_c_20_p N_VDD_c_58_n 3.86251e-19
cc_21 N_VSS_c_4_p N_VDD_c_60_n 0.00116512f
cc_22 N_VSS_c_6_p N_VDD_c_61_n 3.44698e-19
cc_23 N_VSS_c_13_p N_VDD_c_61_n 6.36088e-19
cc_24 N_VSS_c_6_p N_B_c_85_n 2.00737e-19
cc_25 N_VSS_c_13_p N_B_c_85_n 2.34295e-19
cc_26 N_VSS_c_4_p N_B_c_85_n 0.0014669f
cc_27 N_VSS_c_6_p N_B_c_88_n 2.15082e-19
cc_28 N_VSS_c_13_p N_B_c_88_n 5.20396e-19
cc_29 N_VSS_c_8_p N_Z_c_105_n 3.43419e-19
cc_30 N_VSS_c_3_p N_Z_c_105_n 3.48267e-19
cc_31 N_VSS_c_31_p N_Z_c_107_n 3.43419e-19
cc_32 N_VSS_c_32_p N_Z_c_107_n 3.48267e-19
cc_33 N_VSS_c_8_p N_Z_c_109_n 3.48267e-19
cc_34 N_VSS_c_31_p N_Z_c_109_n 3.48267e-19
cc_35 N_VSS_c_3_p N_Z_c_109_n 8.54909e-19
cc_36 N_VSS_c_32_p N_Z_c_109_n 5.71987e-19
cc_37 N_VSS_c_4_p N_Z_c_109_n 0.00105386f
cc_38 N_VSS_c_15_p N_Z_c_109_n 2.24858e-19
cc_39 N_VSS_XI6.X0_PGD N_A_c_129_n 7.89465e-19
cc_40 N_VDD_c_63_p N_B_c_90_n 4.99294e-19
cc_41 N_VDD_c_42_n N_B_c_85_n 0.0026351f
cc_42 N_VDD_c_65_p N_B_c_85_n 3.50338e-19
cc_43 N_VDD_c_66_p N_B_c_85_n 2.36346e-19
cc_44 N_VDD_c_42_n N_B_c_94_n 5.07158e-19
cc_45 N_VDD_c_65_p N_B_c_94_n 2.30903e-19
cc_46 N_VDD_c_42_n N_B_c_88_n 3.66936e-19
cc_47 N_VDD_c_70_p N_Z_c_107_n 3.43419e-19
cc_48 N_VDD_c_49_n N_Z_c_107_n 3.72199e-19
cc_49 N_VDD_c_50_n N_Z_c_107_n 2.74986e-19
cc_50 N_VDD_c_70_p N_Z_c_109_n 3.48267e-19
cc_51 N_VDD_c_42_n N_Z_c_109_n 0.00130587f
cc_52 N_VDD_c_49_n N_Z_c_109_n 7.92786e-19
cc_53 N_VDD_c_50_n N_Z_c_109_n 3.84599e-19
cc_54 N_VDD_XI8.X0_PGD N_A_c_129_n 5.98669e-19
cc_55 N_VDD_XI7.X0_PGD N_A_c_129_n 2.07763e-19
cc_56 N_VDD_XI8.X0_PGS N_A_c_132_n 8.07534e-19
cc_57 N_VDD_c_42_n N_A_c_132_n 5.64288e-19
cc_58 N_VDD_c_58_n N_A_c_134_n 2.30699e-19
cc_59 N_VDD_c_61_n N_A_c_134_n 5.11881e-19
cc_60 N_VDD_c_58_n N_A_c_136_n 2.87155e-19
cc_61 N_VDD_c_61_n N_A_c_136_n 2.16965e-19
cc_62 N_B_c_85_n N_Z_c_109_n 0.00740143f
cc_63 N_B_c_94_n N_Z_c_109_n 0.0010409f
cc_64 N_B_c_88_n N_Z_c_109_n 9.58642e-19
cc_65 N_B_c_100_p N_A_XI6.X0_PGS 4.87172e-19
cc_66 N_B_c_88_n N_A_XI6.X0_PGS 0.00109812f
cc_67 N_B_c_94_n N_A_c_129_n 0.00222679f
cc_68 N_B_c_88_n N_A_c_129_n 4.51405e-19
cc_69 N_B_c_88_n N_A_c_134_n 8.88364e-19
cc_70 N_Z_c_107_n N_A_c_129_n 4.45349e-19
cc_71 N_Z_c_109_n N_A_c_129_n 9.69188e-19
cc_72 N_Z_c_109_n N_A_c_134_n 0.00114087f
cc_73 N_Z_c_109_n N_A_c_136_n 0.00155484f
*
.ends
*
*
.subckt NOR2_HPNW12 A B Y VDD VSS
xgate (VSS VDD B Y A) G2_NOR2_N3
.ends
*
* File: G2_OAI21_N3.pex.netlist
* Created: Wed Mar  2 11:39:40 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_OAI21_N3_VSS 2 4 6 8 10 22 29 37 42 45 50 55 64 73 74 78 84 86 91
+ 94 Vss
c48 92 Vss 5.73928e-19
c49 91 Vss 0.00930467f
c50 86 Vss 0.00178323f
c51 84 Vss 0.00287693f
c52 79 Vss 0.00137325f
c53 78 Vss 0.00727688f
c54 74 Vss 6.08576e-19
c55 73 Vss 0.00762928f
c56 64 Vss 0.00685524f
c57 55 Vss 2.01979e-19
c58 50 Vss 0.00208662f
c59 45 Vss 0.00137663f
c60 42 Vss 0.00818763f
c61 37 Vss 0.00963114f
c62 33 Vss 0.0307825f
c63 29 Vss 5.22622e-20
c64 26 Vss 0.101261f
c65 22 Vss 0.0345879f
c66 21 Vss 0.0712517f
c67 10 Vss 0.191158f
c68 8 Vss 0.19018f
c69 4 Vss 0.189789f
r70 91 94 0.326018
r71 90 91 18.8387
r72 86 90 0.655813
r73 85 92 0.494161
r74 84 94 0.326018
r75 84 85 4.33457
r76 80 92 0.128424
r77 78 92 0.494161
r78 78 79 10.1696
r79 73 79 0.652036
r80 72 74 0.655813
r81 72 73 18.8387
r82 55 86 1.82344
r83 50 64 1.16709
r84 50 80 2.16729
r85 45 74 1.82344
r86 42 55 1.16709
r87 37 45 1.16709
r88 29 64 0.238214
r89 27 33 0.494161
r90 27 29 1.5171
r91 26 30 0.652036
r92 26 29 1.4004
r93 23 33 0.128424
r94 21 33 0.494161
r95 21 22 2.8008
r96 18 22 0.652036
r97 10 30 5.1348
r98 8 23 5.1348
r99 6 42 0.123773
r100 4 18 5.1348
r101 2 37 0.123773
.ends

.subckt PM_G2_OAI21_N3_VDD 2 4 6 8 30 35 38 39 41 43 49 51 56 59 65 Vss
c48 65 Vss 0.00671256f
c49 57 Vss 5.35171e-19
c50 56 Vss 0.0125966f
c51 55 Vss 0.0017875f
c52 51 Vss 0.00240793f
c53 49 Vss 0.00382188f
c54 47 Vss 0.00183797f
c55 43 Vss 0.00172744f
c56 41 Vss 8.2329e-19
c57 40 Vss 0.0017875f
c58 39 Vss 0.00981811f
c59 38 Vss 0.0129397f
c60 35 Vss 0.00815963f
c61 30 Vss 0.0082356f
c62 25 Vss 0.0855608f
c63 19 Vss 0.034095f
c64 18 Vss 0.0688526f
c65 6 Vss 0.192138f
c66 2 Vss 0.192543f
r67 55 59 0.326018
r68 55 56 18.8804
r69 51 56 0.655813
r70 51 53 1.82344
r71 50 57 0.494161
r72 49 59 0.326018
r73 49 50 4.37625
r74 47 65 1.16709
r75 45 57 0.128424
r76 45 47 2.20896
r77 41 43 1.82344
r78 39 57 0.494161
r79 39 40 10.1279
r80 38 41 0.655813
r81 37 40 0.652036
r82 37 38 18.8804
r83 35 53 1.16709
r84 30 43 1.16709
r85 25 65 0.238214
r86 23 25 2.04225
r87 20 23 0.0685365
r88 18 23 0.5835
r89 18 19 2.8008
r90 15 19 0.652036
r91 8 35 0.123773
r92 6 20 5.1348
r93 4 30 0.123773
r94 2 15 5.1348
.ends

.subckt PM_G2_OAI21_N3_B 2 4 13 18 21 26 31 Vss
c19 31 Vss 0.00415668f
c20 26 Vss 0.0032846f
c21 18 Vss 9.6577e-19
c22 13 Vss 0.167996f
c23 2 Vss 0.166757f
r24 23 31 1.16709
r25 21 23 1.66714
r26 18 26 1.16709
r27 18 21 3.16757
r28 13 31 0.476429
r29 10 26 0.50025
r30 4 13 4.4346
r31 2 10 4.37625
.ends

.subckt PM_G2_OAI21_N3_A 2 4 13 18 21 26 31 36 44 46 Vss
c38 46 Vss 1.44014e-19
c39 36 Vss 0.00294987f
c40 31 Vss 0.00806931f
c41 26 Vss 0.0038514f
c42 21 Vss 0.00314266f
c43 18 Vss 0.0859029f
c44 13 Vss 4.64808e-20
c45 4 Vss 0.166608f
c46 2 Vss 0.193159f
r47 40 46 0.655813
r48 26 36 1.16709
r49 26 46 4.52212
r50 21 31 1.16709
r51 21 44 0.0833571
r52 21 40 12.6703
r53 18 31 0.238214
r54 15 18 1.92555
r55 13 36 0.50025
r56 7 15 0.0685365
r57 4 13 4.37625
r58 2 7 5.1348
.ends

.subckt PM_G2_OAI21_N3_Z 2 4 6 8 23 27 30 33 Vss
c33 30 Vss 0.0016158f
c34 27 Vss 0.00640524f
c35 23 Vss 0.00630974f
c36 8 Vss 0.00143493f
c37 6 Vss 0.00143493f
r38 33 35 7.54382
r39 30 33 5.29318
r40 27 35 1.16709
r41 23 30 1.16709
r42 8 27 0.123773
r43 6 23 0.123773
r44 4 27 0.123773
r45 2 23 0.123773
.ends

.subckt PM_G2_OAI21_N3_C 2 4 6 13 14 17 24 27 Vss
c28 27 Vss 7.80628e-19
c29 24 Vss 0.0813012f
c30 17 Vss 0.25734f
c31 14 Vss 0.0348849f
c32 13 Vss 0.247183f
c33 4 Vss 0.29011f
c34 2 Vss 0.290309f
r35 27 30 0.0833571
r36 23 24 2.04225
r37 20 24 0.0685365
r38 17 30 1.16709
r39 15 23 0.0685365
r40 15 17 2.8008
r41 13 23 0.5835
r42 13 14 8.92755
r43 10 14 0.652036
r44 6 17 5.6016
r45 4 20 8.4024
r46 2 10 8.4024
.ends

.subckt G2_OAI21_N3  VSS VDD B A Z C
*
* C	C
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI7.X0 N_Z_XI7.X0_D N_VDD_XI7.X0_PGD N_B_XI7.X0_CG N_C_XI7.X0_PGS N_VSS_XI7.X0_S
+ TIGFET_HPNW12
XI5.X0 N_Z_XI5.X0_D N_VSS_XI5.X0_PGD N_B_XI5.X0_CG N_A_XI5.X0_PGS N_VDD_XI5.X0_S
+ TIGFET_HPNW12
XI8.X0 N_Z_XI8.X0_D N_VDD_XI8.X0_PGD N_A_XI8.X0_CG N_C_XI8.X0_PGS N_VSS_XI8.X0_S
+ TIGFET_HPNW12
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_C_XI6.X0_CG N_VSS_XI6.X0_PGS
+ N_VDD_XI6.X0_S TIGFET_HPNW12
*
x_PM_G2_OAI21_N3_VSS N_VSS_XI7.X0_S N_VSS_XI5.X0_PGD N_VSS_XI8.X0_S
+ N_VSS_XI6.X0_PGD N_VSS_XI6.X0_PGS N_VSS_c_30_p N_VSS_c_46_p N_VSS_c_1_p
+ N_VSS_c_10_p N_VSS_c_2_p N_VSS_c_22_p N_VSS_c_11_p N_VSS_c_23_p N_VSS_c_3_p
+ N_VSS_c_4_p N_VSS_c_9_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_15_p VSS Vss
+ PM_G2_OAI21_N3_VSS
x_PM_G2_OAI21_N3_VDD N_VDD_XI7.X0_PGD N_VDD_XI5.X0_S N_VDD_XI8.X0_PGD
+ N_VDD_XI6.X0_S N_VDD_c_80_p N_VDD_c_81_p N_VDD_c_49_n N_VDD_c_53_n
+ N_VDD_c_55_n N_VDD_c_56_n N_VDD_c_58_n N_VDD_c_61_n N_VDD_c_64_n VDD
+ N_VDD_c_71_p Vss PM_G2_OAI21_N3_VDD
x_PM_G2_OAI21_N3_B N_B_XI7.X0_CG N_B_XI5.X0_CG N_B_c_103_p N_B_c_97_n B
+ N_B_c_99_n N_B_c_100_n Vss PM_G2_OAI21_N3_B
x_PM_G2_OAI21_N3_A N_A_XI5.X0_PGS N_A_XI8.X0_CG N_A_c_130_n N_A_c_137_n
+ N_A_c_117_n N_A_c_122_n N_A_c_124_n N_A_c_134_n A N_A_c_128_n Vss
+ PM_G2_OAI21_N3_A
x_PM_G2_OAI21_N3_Z N_Z_XI7.X0_D N_Z_XI5.X0_D N_Z_XI8.X0_D N_Z_XI6.X0_D
+ N_Z_c_154_n N_Z_c_165_n N_Z_c_158_n Z Vss PM_G2_OAI21_N3_Z
x_PM_G2_OAI21_N3_C N_C_XI7.X0_PGS N_C_XI8.X0_PGS N_C_XI6.X0_CG N_C_c_187_n
+ N_C_c_206_n N_C_c_189_n N_C_c_191_n C Vss PM_G2_OAI21_N3_C
cc_1 N_VSS_c_1_p N_VDD_c_49_n 9.5668e-19
cc_2 N_VSS_c_2_p N_VDD_c_49_n 0.00165395f
cc_3 N_VSS_c_3_p N_VDD_c_49_n 0.00820308f
cc_4 N_VSS_c_4_p N_VDD_c_49_n 0.00189979f
cc_5 N_VSS_c_1_p N_VDD_c_53_n 2.43883e-19
cc_6 N_VSS_c_2_p N_VDD_c_53_n 7.51487e-19
cc_7 N_VSS_c_3_p N_VDD_c_55_n 0.00170274f
cc_8 N_VSS_c_2_p N_VDD_c_56_n 4.01889e-19
cc_9 N_VSS_c_9_p N_VDD_c_56_n 4.74109e-19
cc_10 N_VSS_c_10_p N_VDD_c_58_n 2.43883e-19
cc_11 N_VSS_c_11_p N_VDD_c_58_n 3.33988e-19
cc_12 N_VSS_c_12_p N_VDD_c_58_n 4.17499e-19
cc_13 N_VSS_c_13_p N_VDD_c_61_n 4.74109e-19
cc_14 N_VSS_c_12_p N_VDD_c_61_n 4.01889e-19
cc_15 N_VSS_c_15_p N_VDD_c_61_n 0.00178085f
cc_16 N_VSS_c_10_p N_VDD_c_64_n 9.5668e-19
cc_17 N_VSS_c_11_p N_VDD_c_64_n 0.00165395f
cc_18 N_VSS_c_12_p N_VDD_c_64_n 0.00189979f
cc_19 N_VSS_c_15_p N_VDD_c_64_n 0.0087982f
cc_20 N_VSS_c_3_p N_B_c_97_n 5.69535e-19
cc_21 N_VSS_XI5.X0_PGD N_A_XI5.X0_PGS 0.00176902f
cc_22 N_VSS_c_22_p N_A_c_117_n 8.59446e-19
cc_23 N_VSS_c_23_p N_A_c_117_n 3.44698e-19
cc_24 N_VSS_c_3_p N_A_c_117_n 0.00485346f
cc_25 N_VSS_c_9_p N_A_c_117_n 0.00211426f
cc_26 N_VSS_c_15_p N_A_c_117_n 0.00226606f
cc_27 N_VSS_c_9_p N_A_c_122_n 6.38907e-19
cc_28 N_VSS_c_15_p N_A_c_122_n 7.9739e-19
cc_29 N_VSS_XI5.X0_PGD N_A_c_124_n 3.11814e-19
cc_30 N_VSS_c_30_p N_A_c_124_n 0.00322564f
cc_31 N_VSS_c_22_p N_A_c_124_n 3.44698e-19
cc_32 N_VSS_c_23_p N_A_c_124_n 6.61253e-19
cc_33 N_VSS_c_3_p N_A_c_128_n 0.00309992f
cc_34 N_VSS_c_1_p N_Z_c_154_n 3.43419e-19
cc_35 N_VSS_c_10_p N_Z_c_154_n 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_c_154_n 3.48267e-19
cc_37 N_VSS_c_11_p N_Z_c_154_n 3.48267e-19
cc_38 N_VSS_c_1_p N_Z_c_158_n 3.48267e-19
cc_39 N_VSS_c_10_p N_Z_c_158_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_158_n 5.71987e-19
cc_41 N_VSS_c_11_p N_Z_c_158_n 5.71987e-19
cc_42 N_VSS_c_9_p N_Z_c_158_n 3.21537e-19
cc_43 N_VSS_c_15_p N_Z_c_158_n 8.14216e-19
cc_44 N_VSS_XI5.X0_PGD N_C_c_187_n 6.83817e-19
cc_45 N_VSS_XI6.X0_PGD N_C_c_187_n 6.83817e-19
cc_46 N_VSS_c_46_p N_C_c_189_n 2.53848e-19
cc_47 N_VSS_c_23_p N_C_c_189_n 0.00232974f
cc_48 N_VSS_XI6.X0_PGS N_C_c_191_n 8.42974e-19
cc_49 N_VDD_c_49_n N_B_c_97_n 0.00231792f
cc_50 N_VDD_c_49_n N_B_c_99_n 3.66936e-19
cc_51 N_VDD_c_49_n N_B_c_100_n 4.8547e-19
cc_52 N_VDD_c_71_p N_A_XI8.X0_CG 0.00266603f
cc_53 N_VDD_c_71_p N_A_c_130_n 5.2106e-19
cc_54 N_VDD_c_53_n N_A_c_122_n 6.20865e-19
cc_55 N_VDD_c_64_n N_A_c_122_n 6.23587e-19
cc_56 N_VDD_c_71_p N_A_c_122_n 2.23358e-19
cc_57 N_VDD_c_64_n N_A_c_134_n 3.66936e-19
cc_58 N_VDD_c_71_p N_A_c_134_n 3.65437e-19
cc_59 N_VDD_c_49_n N_A_c_128_n 6.11072e-19
cc_60 N_VDD_c_53_n N_Z_c_154_n 2.43883e-19
cc_61 N_VDD_c_80_p N_Z_c_165_n 3.43419e-19
cc_62 N_VDD_c_81_p N_Z_c_165_n 3.43419e-19
cc_63 N_VDD_c_56_n N_Z_c_165_n 3.72199e-19
cc_64 N_VDD_c_61_n N_Z_c_165_n 3.72199e-19
cc_65 N_VDD_c_80_p N_Z_c_158_n 3.48267e-19
cc_66 N_VDD_c_81_p N_Z_c_158_n 3.48267e-19
cc_67 N_VDD_c_49_n N_Z_c_158_n 0.00116129f
cc_68 N_VDD_c_53_n N_Z_c_158_n 5.05821e-19
cc_69 N_VDD_c_56_n N_Z_c_158_n 5.09542e-19
cc_70 N_VDD_c_61_n N_Z_c_158_n 7.72285e-19
cc_71 N_VDD_c_64_n N_Z_c_158_n 0.00182594f
cc_72 N_VDD_c_49_n N_C_XI7.X0_PGS 6.13097e-19
cc_73 N_VDD_c_64_n N_C_XI8.X0_PGS 6.32546e-19
cc_74 N_VDD_XI7.X0_PGD N_C_c_187_n 6.83817e-19
cc_75 N_VDD_XI8.X0_PGD N_C_c_187_n 6.83817e-19
cc_76 N_VDD_c_64_n N_C_c_189_n 5.92666e-19
cc_77 N_VDD_c_64_n C 5.04211e-19
cc_78 N_B_c_100_n N_A_c_137_n 2.60115e-19
cc_79 N_B_c_97_n N_A_c_117_n 0.00265561f
cc_80 N_B_c_103_p N_A_c_124_n 0.00262973f
cc_81 N_B_c_97_n N_A_c_124_n 2.40146e-19
cc_82 N_B_c_100_n N_A_c_124_n 3.65437e-19
cc_83 N_B_c_99_n N_A_c_134_n 8.86454e-19
cc_84 N_B_c_97_n N_A_c_128_n 7.49556e-19
cc_85 N_B_c_97_n N_Z_c_158_n 0.00671f
cc_86 N_B_c_99_n N_Z_c_158_n 9.58174e-19
cc_87 N_B_c_100_n N_Z_c_158_n 0.00101748f
cc_88 N_B_XI7.X0_CG N_C_XI7.X0_PGS 4.87172e-19
cc_89 N_B_c_99_n N_C_XI7.X0_PGS 0.001089f
cc_90 N_B_c_99_n N_C_c_187_n 6.02551e-19
cc_91 N_B_c_100_n N_C_c_187_n 0.00149356f
cc_92 N_B_c_100_n N_C_c_189_n 9.54365e-19
cc_93 N_A_c_117_n N_Z_c_158_n 0.00195546f
cc_94 N_A_c_122_n N_Z_c_158_n 0.00358051f
cc_95 N_A_c_134_n N_Z_c_158_n 9.53427e-19
cc_96 N_A_XI8.X0_CG N_C_XI8.X0_PGS 4.87172e-19
cc_97 N_A_c_134_n N_C_XI8.X0_PGS 0.001089f
cc_98 N_A_c_134_n N_C_c_187_n 0.00157146f
cc_99 N_A_XI5.X0_PGS N_C_c_206_n 8.42974e-19
cc_100 N_A_c_122_n N_C_c_189_n 5.38228e-19
cc_101 N_A_c_134_n N_C_c_189_n 0.00222154f
cc_102 N_A_c_122_n C 8.18489e-19
cc_103 N_Z_c_154_n N_C_c_187_n 3.5202e-19
cc_104 N_Z_c_165_n N_C_c_187_n 3.5202e-19
cc_105 N_Z_c_158_n N_C_c_187_n 3.56555e-19
cc_106 N_Z_c_158_n N_C_c_189_n 0.00101565f
cc_107 N_Z_c_158_n C 0.00141616f
*
.ends
*
*
.subckt OAI21_HPNW12 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 A0 Y B0) G2_OAI21_N3
.ends
*
* File: G3_OR2_N3.pex.netlist
* Created: Tue Mar  1 12:18:46 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_OR2_N3_VSS 2 4 6 8 10 12 28 29 38 44 49 52 57 62 67 76 85 90 91 95
+ 96 101 107 114 115 116 Vss
c71 116 Vss 3.91906e-19
c72 115 Vss 3.75522e-19
c73 107 Vss 0.00372185f
c74 101 Vss 0.00290457f
c75 96 Vss 8.35017e-19
c76 95 Vss 0.00178035f
c77 91 Vss 6.20207e-19
c78 90 Vss 0.00579798f
c79 85 Vss 0.0039758f
c80 76 Vss 0.0050462f
c81 67 Vss 5.89061e-19
c82 62 Vss 8.97934e-19
c83 57 Vss 0.00103095f
c84 52 Vss 0.00124124f
c85 49 Vss 0.00687623f
c86 44 Vss 0.00812495f
c87 38 Vss 0.0895788f
c88 29 Vss 0.0349332f
c89 28 Vss 0.0997249f
c90 12 Vss 0.190073f
c91 10 Vss 0.189045f
c92 8 Vss 0.00143493f
c93 4 Vss 0.189407f
r94 109 114 0.458464
r95 108 116 0.494161
r96 107 109 0.652036
r97 107 108 7.46046
r98 103 116 0.128424
r99 102 115 0.494161
r100 101 116 0.494161
r101 101 102 7.46046
r102 97 115 0.128424
r103 95 115 0.494161
r104 95 96 4.37625
r105 90 96 0.652036
r106 89 91 0.655813
r107 89 90 18.3386
r108 67 85 1.16709
r109 67 114 1.70882
r110 62 103 6.16843
r111 57 76 1.16709
r112 57 97 2.16729
r113 52 91 1.82344
r114 49 62 1.16709
r115 44 52 1.16709
r116 36 76 0.0476429
r117 36 38 2.04225
r118 31 85 0.0476429
r119 29 31 1.45875
r120 28 32 0.652036
r121 28 31 1.45875
r122 25 29 0.652036
r123 22 38 0.0685365
r124 12 32 5.1348
r125 10 25 5.1348
r126 8 49 0.123773
r127 6 49 0.123773
r128 4 22 5.1348
r129 2 44 0.123773
.ends

.subckt PM_G3_OR2_N3_VDD 2 4 6 8 10 12 14 16 37 46 56 62 67 70 72 73 77 79 80 83
+ 87 89 93 95 97 102 103 104 105 107 113 119 124 Vss
c78 124 Vss 0.00450608f
c79 119 Vss 0.00587228f
c80 113 Vss 0.00493107f
c81 105 Vss 2.39889e-19
c82 104 Vss 2.39889e-19
c83 103 Vss 4.52364e-19
c84 102 Vss 0.00430335f
c85 101 Vss 0.00170674f
c86 97 Vss 0.00160078f
c87 95 Vss 0.00854117f
c88 93 Vss 7.28478e-19
c89 89 Vss 0.00205766f
c90 87 Vss 4.80319e-19
c91 83 Vss 0.00133062f
c92 80 Vss 8.68835e-19
c93 79 Vss 0.00561215f
c94 77 Vss 0.0017471f
c95 74 Vss 0.00174847f
c96 73 Vss 0.00498635f
c97 72 Vss 0.00313638f
c98 70 Vss 0.0119561f
c99 67 Vss 0.0100342f
c100 62 Vss 0.00818522f
c101 57 Vss 0.129193f
c102 56 Vss 7.73513e-20
c103 47 Vss 0.035874f
c104 46 Vss 0.101312f
c105 37 Vss 0.0356247f
c106 36 Vss 0.101564f
c107 14 Vss 0.189069f
c108 12 Vss 0.189513f
c109 10 Vss 0.189312f
c110 8 Vss 0.189362f
c111 4 Vss 0.191197f
c112 2 Vss 0.192293f
r113 113 116 0.05
r114 101 107 0.349767
r115 101 102 5.50157
r116 97 107 0.306046
r117 97 99 1.82344
r118 96 105 0.494161
r119 95 102 0.652036
r120 95 96 10.1279
r121 93 124 1.16709
r122 91 105 0.128424
r123 91 93 2.16729
r124 90 104 0.494161
r125 89 105 0.494161
r126 89 90 4.54296
r127 87 119 1.16709
r128 85 104 0.128424
r129 85 87 2.16729
r130 83 116 1.16709
r131 81 83 2.16729
r132 79 104 0.494161
r133 79 80 10.1696
r134 75 103 0.0828784
r135 75 77 1.82344
r136 73 81 0.652036
r137 73 74 4.37625
r138 72 80 0.652036
r139 71 103 0.551426
r140 71 72 5.50157
r141 70 103 0.551426
r142 69 74 0.652036
r143 69 70 18.2969
r144 67 99 1.16709
r145 62 77 1.16709
r146 56 113 0.0238214
r147 56 57 2.26917
r148 53 56 2.26917
r149 49 124 0.0476429
r150 47 49 1.45875
r151 46 50 0.652036
r152 46 49 1.45875
r153 43 47 0.652036
r154 39 119 0.0476429
r155 37 39 1.5171
r156 36 40 0.652036
r157 36 39 1.4004
r158 33 37 0.652036
r159 30 57 0.00605528
r160 27 53 0.00605528
r161 16 67 0.123773
r162 14 43 5.1348
r163 12 50 5.1348
r164 10 40 5.1348
r165 8 33 5.1348
r166 6 62 0.123773
r167 4 27 5.1348
r168 2 30 5.1348
.ends

.subckt PM_G3_OR2_N3_B 2 4 10 13 18 21 26 31 Vss
c19 31 Vss 0.00192399f
c20 26 Vss 0.00378619f
c21 18 Vss 0.00125219f
c22 13 Vss 0.166574f
c23 10 Vss 7.84101e-20
c24 2 Vss 0.16675f
r25 23 31 1.16709
r26 21 23 2.29232
r27 18 26 1.16709
r28 18 21 2.54239
r29 13 31 0.50025
r30 10 26 0.50025
r31 4 13 4.37625
r32 2 10 4.37625
.ends

.subckt PM_G3_OR2_N3_NET21 2 4 6 8 10 24 27 38 42 45 53 66 70 Vss
c35 70 Vss 0.00748471f
c36 66 Vss 0.00592889f
c37 53 Vss 0.0020112f
c38 45 Vss 0.00308864f
c39 42 Vss 0.00545637f
c40 38 Vss 0.00813452f
c41 27 Vss 8.95828e-20
c42 24 Vss 0.229828f
c43 21 Vss 0.18045f
c44 19 Vss 0.0247918f
c45 10 Vss 0.193588f
c46 6 Vss 0.00143493f
r47 70 74 0.652036
r48 53 66 1.16709
r49 53 74 2.16729
r50 48 70 8.04396
r51 48 50 6.75193
r52 45 48 6.08507
r53 42 50 1.16709
r54 38 45 1.16709
r55 27 66 0.0476429
r56 25 27 0.326018
r57 25 27 0.1167
r58 24 28 0.652036
r59 24 27 6.7686
r60 21 66 0.357321
r61 19 27 0.326018
r62 19 21 0.40845
r63 10 28 5.1348
r64 8 21 4.72635
r65 6 42 0.123773
r66 4 42 0.123773
r67 2 38 0.123773
.ends

.subckt PM_G3_OR2_N3_A 2 4 10 11 14 18 21 Vss
c21 18 Vss 3.08468e-19
c22 14 Vss 0.225307f
c23 11 Vss 0.0348763f
c24 10 Vss 0.278488f
c25 2 Vss 0.253009f
r26 18 27 1.16709
r27 18 21 0.0416786
r28 14 27 0.05
r29 12 14 1.6338
r30 10 12 0.652036
r31 10 11 8.92755
r32 7 11 0.652036
r33 4 14 5.6016
r34 2 7 7.2354
.ends

.subckt PM_G3_OR2_N3_Z 2 4 13 19 Vss
c12 13 Vss 0.00498872f
c13 4 Vss 0.00143493f
r14 16 19 0.0364688
r15 13 16 1.16709
r16 4 13 0.123773
r17 2 13 0.123773
.ends

.subckt G3_OR2_N3  VSS VDD B A Z
*
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI12.X0 N_NET21_XI12.X0_D N_VDD_XI12.X0_PGD N_B_XI12.X0_CG N_VDD_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW12
XI10.X0 N_NET21_XI10.X0_D N_VSS_XI10.X0_PGD N_B_XI10.X0_CG N_A_XI10.X0_PGS
+ N_VDD_XI10.X0_S TIGFET_HPNW12
XI11.X0 N_NET21_XI11.X0_D N_VDD_XI11.X0_PGD N_A_XI11.X0_CG N_VDD_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW12
XI14.X0 N_Z_XI14.X0_D N_VDD_XI14.X0_PGD N_NET21_XI14.X0_CG N_VDD_XI14.X0_PGS
+ N_VSS_XI14.X0_S TIGFET_HPNW12
XI13.X0 N_Z_XI13.X0_D N_VSS_XI13.X0_PGD N_NET21_XI13.X0_CG N_VSS_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW12
*
x_PM_G3_OR2_N3_VSS N_VSS_XI12.X0_S N_VSS_XI10.X0_PGD N_VSS_XI11.X0_S
+ N_VSS_XI14.X0_S N_VSS_XI13.X0_PGD N_VSS_XI13.X0_PGS N_VSS_c_32_p N_VSS_c_4_p
+ N_VSS_c_3_p N_VSS_c_11_p N_VSS_c_24_p N_VSS_c_5_p N_VSS_c_8_p N_VSS_c_22_p
+ N_VSS_c_30_p N_VSS_c_9_p N_VSS_c_31_p N_VSS_c_6_p N_VSS_c_7_p N_VSS_c_17_p
+ N_VSS_c_20_p N_VSS_c_18_p N_VSS_c_27_p VSS N_VSS_c_19_p N_VSS_c_28_p Vss
+ PM_G3_OR2_N3_VSS
x_PM_G3_OR2_N3_VDD N_VDD_XI12.X0_PGD N_VDD_XI12.X0_PGS N_VDD_XI10.X0_S
+ N_VDD_XI11.X0_PGD N_VDD_XI11.X0_PGS N_VDD_XI14.X0_PGD N_VDD_XI14.X0_PGS
+ N_VDD_XI13.X0_S N_VDD_c_74_n N_VDD_c_75_n N_VDD_c_119_p N_VDD_c_128_p
+ N_VDD_c_144_p N_VDD_c_76_n N_VDD_c_79_n N_VDD_c_82_n N_VDD_c_84_n N_VDD_c_85_n
+ N_VDD_c_91_n N_VDD_c_121_p N_VDD_c_92_n N_VDD_c_95_n N_VDD_c_100_n
+ N_VDD_c_103_n N_VDD_c_146_p N_VDD_c_108_n N_VDD_c_112_n N_VDD_c_113_n
+ N_VDD_c_114_n VDD N_VDD_c_122_p N_VDD_c_115_n N_VDD_c_117_n Vss
+ PM_G3_OR2_N3_VDD
x_PM_G3_OR2_N3_B N_B_XI12.X0_CG N_B_XI10.X0_CG N_B_c_155_n N_B_c_165_p
+ N_B_c_150_n B N_B_c_159_n N_B_c_153_n Vss PM_G3_OR2_N3_B
x_PM_G3_OR2_N3_NET21 N_NET21_XI12.X0_D N_NET21_XI10.X0_D N_NET21_XI11.X0_D
+ N_NET21_XI14.X0_CG N_NET21_XI13.X0_CG N_NET21_c_169_n N_NET21_c_183_n
+ N_NET21_c_170_n N_NET21_c_172_n N_NET21_c_174_n N_NET21_c_191_n
+ N_NET21_c_199_p N_NET21_c_179_n Vss PM_G3_OR2_N3_NET21
x_PM_G3_OR2_N3_A N_A_XI10.X0_PGS N_A_XI11.X0_CG N_A_c_204_n N_A_c_207_n
+ N_A_c_209_n N_A_c_211_n A Vss PM_G3_OR2_N3_A
x_PM_G3_OR2_N3_Z N_Z_XI14.X0_D N_Z_XI13.X0_D N_Z_c_225_n Z Vss PM_G3_OR2_N3_Z
cc_1 N_VSS_XI10.X0_PGD N_VDD_XI11.X0_PGD 0.00203999f
cc_2 N_VSS_XI13.X0_PGD N_VDD_XI14.X0_PGD 0.00196229f
cc_3 N_VSS_c_3_p N_VDD_c_74_n 0.00203999f
cc_4 N_VSS_c_4_p N_VDD_c_75_n 0.00196229f
cc_5 N_VSS_c_5_p N_VDD_c_76_n 0.00187494f
cc_6 N_VSS_c_6_p N_VDD_c_76_n 0.0079127f
cc_7 N_VSS_c_7_p N_VDD_c_76_n 0.00189882f
cc_8 N_VSS_c_8_p N_VDD_c_79_n 4.35319e-19
cc_9 N_VSS_c_9_p N_VDD_c_79_n 4.7255e-19
cc_10 N_VSS_c_6_p N_VDD_c_79_n 0.00412661f
cc_11 N_VSS_c_11_p N_VDD_c_82_n 2.77593e-19
cc_12 N_VSS_c_5_p N_VDD_c_82_n 8.30039e-19
cc_13 N_VSS_c_5_p N_VDD_c_84_n 4.01154e-19
cc_14 N_VSS_c_3_p N_VDD_c_85_n 3.71132e-19
cc_15 N_VSS_c_8_p N_VDD_c_85_n 0.00141228f
cc_16 N_VSS_c_9_p N_VDD_c_85_n 0.00114511f
cc_17 N_VSS_c_17_p N_VDD_c_85_n 0.00352847f
cc_18 N_VSS_c_18_p N_VDD_c_85_n 0.00442704f
cc_19 N_VSS_c_19_p N_VDD_c_85_n 7.74609e-19
cc_20 N_VSS_c_20_p N_VDD_c_91_n 0.00107113f
cc_21 N_VSS_c_8_p N_VDD_c_92_n 8.39054e-19
cc_22 N_VSS_c_22_p N_VDD_c_92_n 3.93845e-19
cc_23 N_VSS_c_9_p N_VDD_c_92_n 3.95933e-19
cc_24 N_VSS_c_24_p N_VDD_c_95_n 2.74986e-19
cc_25 N_VSS_c_22_p N_VDD_c_95_n 2.9533e-19
cc_26 N_VSS_c_18_p N_VDD_c_95_n 0.00139286f
cc_27 N_VSS_c_27_p N_VDD_c_95_n 0.0014416f
cc_28 N_VSS_c_28_p N_VDD_c_95_n 0.00111918f
cc_29 N_VSS_c_22_p N_VDD_c_100_n 3.91951e-19
cc_30 N_VSS_c_30_p N_VDD_c_100_n 8.45954e-19
cc_31 N_VSS_c_31_p N_VDD_c_100_n 3.99794e-19
cc_32 N_VSS_c_32_p N_VDD_c_103_n 4.0633e-19
cc_33 N_VSS_c_4_p N_VDD_c_103_n 3.89167e-19
cc_34 N_VSS_c_30_p N_VDD_c_103_n 0.00161703f
cc_35 N_VSS_c_31_p N_VDD_c_103_n 2.26455e-19
cc_36 N_VSS_c_27_p N_VDD_c_103_n 0.00619092f
cc_37 N_VSS_XI13.X0_PGS N_VDD_c_108_n 4.28478e-19
cc_38 N_VSS_c_22_p N_VDD_c_108_n 2.85882e-19
cc_39 N_VSS_c_30_p N_VDD_c_108_n 8.67538e-19
cc_40 N_VSS_c_31_p N_VDD_c_108_n 3.66936e-19
cc_41 N_VSS_c_6_p N_VDD_c_112_n 0.00116512f
cc_42 N_VSS_c_18_p N_VDD_c_113_n 0.00102637f
cc_43 N_VSS_c_27_p N_VDD_c_114_n 0.00103008f
cc_44 N_VSS_c_8_p N_VDD_c_115_n 3.44698e-19
cc_45 N_VSS_c_9_p N_VDD_c_115_n 6.36088e-19
cc_46 N_VSS_c_30_p N_VDD_c_117_n 3.48267e-19
cc_47 N_VSS_c_31_p N_VDD_c_117_n 6.489e-19
cc_48 N_VSS_c_8_p N_B_c_150_n 2.0198e-19
cc_49 N_VSS_c_9_p N_B_c_150_n 2.34295e-19
cc_50 N_VSS_c_6_p N_B_c_150_n 9.20502e-19
cc_51 N_VSS_c_8_p N_B_c_153_n 2.15082e-19
cc_52 N_VSS_c_9_p N_B_c_153_n 5.28949e-19
cc_53 N_VSS_XI13.X0_PGD N_NET21_c_169_n 4.31283e-19
cc_54 N_VSS_c_11_p N_NET21_c_170_n 3.43419e-19
cc_55 N_VSS_c_5_p N_NET21_c_170_n 3.48267e-19
cc_56 N_VSS_c_24_p N_NET21_c_172_n 3.43419e-19
cc_57 N_VSS_c_22_p N_NET21_c_172_n 3.48267e-19
cc_58 N_VSS_c_11_p N_NET21_c_174_n 3.48267e-19
cc_59 N_VSS_c_24_p N_NET21_c_174_n 3.48267e-19
cc_60 N_VSS_c_5_p N_NET21_c_174_n 8.54909e-19
cc_61 N_VSS_c_22_p N_NET21_c_174_n 5.71987e-19
cc_62 N_VSS_c_6_p N_NET21_c_174_n 9.99273e-19
cc_63 N_VSS_c_22_p N_NET21_c_179_n 8.10259e-19
cc_64 N_VSS_c_6_p N_NET21_c_179_n 2.03357e-19
cc_65 N_VSS_c_18_p N_NET21_c_179_n 6.96588e-19
cc_66 N_VSS_XI10.X0_PGD N_A_c_204_n 9.58706e-19
cc_67 N_VSS_c_24_p N_Z_c_225_n 3.43419e-19
cc_68 N_VSS_c_22_p N_Z_c_225_n 3.48267e-19
cc_69 N_VSS_c_24_p Z 3.48267e-19
cc_70 N_VSS_c_22_p Z 7.85754e-19
cc_71 N_VSS_c_27_p Z 2.23989e-19
cc_72 N_VDD_c_119_p N_B_c_155_n 5.04908e-19
cc_73 N_VDD_c_76_n N_B_c_150_n 0.00268701f
cc_74 N_VDD_c_121_p N_B_c_150_n 3.49578e-19
cc_75 N_VDD_c_122_p N_B_c_150_n 2.36346e-19
cc_76 N_VDD_c_76_n N_B_c_159_n 5.07158e-19
cc_77 N_VDD_c_121_p N_B_c_159_n 2.30699e-19
cc_78 N_VDD_c_76_n N_B_c_153_n 3.66936e-19
cc_79 N_VDD_XI14.X0_PGD N_NET21_c_169_n 4.31283e-19
cc_80 N_VDD_c_117_n N_NET21_c_183_n 5.33384e-19
cc_81 N_VDD_c_128_p N_NET21_c_172_n 3.43419e-19
cc_82 N_VDD_c_84_n N_NET21_c_172_n 3.72199e-19
cc_83 N_VDD_c_85_n N_NET21_c_172_n 2.74986e-19
cc_84 N_VDD_c_128_p N_NET21_c_174_n 3.48267e-19
cc_85 N_VDD_c_76_n N_NET21_c_174_n 0.00123401f
cc_86 N_VDD_c_84_n N_NET21_c_174_n 7.92786e-19
cc_87 N_VDD_c_85_n N_NET21_c_174_n 3.84599e-19
cc_88 N_VDD_c_117_n N_NET21_c_191_n 2.15082e-19
cc_89 N_VDD_XI12.X0_PGD N_A_c_204_n 5.14897e-19
cc_90 N_VDD_XI11.X0_PGD N_A_c_204_n 2.52296e-19
cc_91 N_VDD_XI12.X0_PGS N_A_c_207_n 6.93093e-19
cc_92 N_VDD_c_76_n N_A_c_207_n 5.08654e-19
cc_93 N_VDD_c_92_n N_A_c_209_n 2.30699e-19
cc_94 N_VDD_c_115_n N_A_c_209_n 5.05291e-19
cc_95 N_VDD_c_92_n N_A_c_211_n 2.64342e-19
cc_96 N_VDD_c_115_n N_A_c_211_n 2.15082e-19
cc_97 N_VDD_c_144_p N_Z_c_225_n 3.43419e-19
cc_98 N_VDD_c_103_n N_Z_c_225_n 2.74986e-19
cc_99 N_VDD_c_146_p N_Z_c_225_n 3.72199e-19
cc_100 N_VDD_c_144_p Z 3.48267e-19
cc_101 N_VDD_c_103_n Z 3.66281e-19
cc_102 N_VDD_c_146_p Z 7.4527e-19
cc_103 N_B_c_150_n N_NET21_c_174_n 0.00754318f
cc_104 N_B_c_159_n N_NET21_c_174_n 0.0010409f
cc_105 N_B_c_153_n N_NET21_c_174_n 9.33005e-19
cc_106 N_B_c_165_p N_A_XI10.X0_PGS 4.87172e-19
cc_107 N_B_c_153_n N_A_XI10.X0_PGS 7.86826e-19
cc_108 N_B_c_159_n N_A_c_204_n 0.00191474f
cc_109 N_B_c_153_n N_A_c_209_n 7.50183e-19
cc_110 N_NET21_c_172_n N_A_c_204_n 4.90018e-19
cc_111 N_NET21_c_174_n N_A_c_204_n 8.56417e-19
cc_112 N_NET21_c_174_n N_A_c_209_n 0.00108943f
cc_113 N_NET21_c_191_n N_A_c_209_n 3.48267e-19
cc_114 N_NET21_c_199_p N_A_c_209_n 0.00171208f
cc_115 N_NET21_c_174_n N_A_c_211_n 0.00142917f
cc_116 N_NET21_c_191_n N_A_c_211_n 4.28721e-19
cc_117 N_NET21_c_179_n N_A_c_211_n 3.71028e-19
cc_118 N_NET21_c_169_n N_Z_c_225_n 7.69306e-19
*
.ends
*
*
.subckt OR2_HPNW12 A B Y VDD VSS
xgate (VSS VDD B A Y) G3_OR2_N3
.ends
*
* File: G4_XNOR2_N3.pex.netlist
* Created: Sun Apr 10 19:31:19 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XNOR2_N3_VDD 2 5 9 12 14 16 32 42 43 45 54 59 66 68 69 70 73 75 76
+ 79 81 85 89 91 93 98 99 100 103 109 114 123 Vss
c102 123 Vss 0.00998345f
c103 114 Vss 0.00466671f
c104 109 Vss 0.00477251f
c105 101 Vss 8.67375e-19
c106 100 Vss 2.39889e-19
c107 99 Vss 4.52364e-19
c108 98 Vss 0.00591503f
c109 93 Vss 0.00301333f
c110 91 Vss 0.0106867f
c111 89 Vss 0.0015063f
c112 85 Vss 6.60056e-19
c113 81 Vss 0.0046084f
c114 79 Vss 0.00109211f
c115 76 Vss 8.68689e-19
c116 75 Vss 0.00224943f
c117 73 Vss 0.00191294f
c118 70 Vss 8.64616e-19
c119 69 Vss 0.00566667f
c120 68 Vss 0.0107726f
c121 66 Vss 0.00280898f
c122 59 Vss 0.00679236f
c123 54 Vss 0.010135f
c124 45 Vss 1.08186e-19
c125 43 Vss 0.0351405f
c126 42 Vss 0.100973f
c127 33 Vss 0.0359366f
c128 32 Vss 0.100971f
c129 14 Vss 0.00143493f
c130 9 Vss 0.377348f
c131 5 Vss 0.379154f
r132 98 103 0.326018
r133 97 98 5.54325
r134 95 123 1.16709
r135 93 97 0.655813
r136 93 95 1.82344
r137 92 101 0.494161
r138 91 103 0.326018
r139 91 92 13.0037
r140 87 101 0.128424
r141 87 89 6.16843
r142 85 114 1.16709
r143 83 85 2.16729
r144 82 100 0.494161
r145 81 101 0.494161
r146 81 82 7.46046
r147 79 109 1.16709
r148 77 100 0.128424
r149 77 79 2.16729
r150 75 100 0.494161
r151 75 76 4.37625
r152 71 99 0.0828784
r153 71 73 1.82344
r154 69 83 0.652036
r155 69 70 10.1279
r156 68 76 0.652036
r157 67 99 0.551426
r158 67 68 17.4633
r159 66 99 0.551426
r160 65 70 0.652036
r161 65 66 5.50157
r162 63 123 0.05
r163 59 89 1.16709
r164 54 73 1.16709
r165 45 114 0.0476429
r166 43 45 1.45875
r167 42 46 0.652036
r168 42 45 1.45875
r169 39 43 0.652036
r170 35 109 0.0476429
r171 33 35 1.45875
r172 32 36 0.652036
r173 32 35 1.45875
r174 29 33 0.652036
r175 16 63 0.123773
r176 14 59 0.123773
r177 12 59 0.123773
r178 9 46 5.1348
r179 9 39 5.1348
r180 5 36 5.1348
r181 5 29 5.1348
r182 2 54 0.123773
.ends

.subckt PM_G4_XNOR2_N3_VSS 3 6 8 11 14 16 32 33 42 43 54 59 63 66 71 76 81 87 96
+ 101 114 116 117 118 123 124 129 137 142 143 144 146 Vss
c85 144 Vss 3.75522e-19
c86 143 Vss 4.28045e-19
c87 142 Vss 0.0047306f
c88 137 Vss 0.00122865f
c89 129 Vss 0.0130341f
c90 124 Vss 8.2479e-19
c91 123 Vss 0.00464476f
c92 118 Vss 8.46757e-19
c93 117 Vss 0.00174235f
c94 116 Vss 0.00202335f
c95 114 Vss 0.00643502f
c96 101 Vss 0.00391102f
c97 96 Vss 0.00421609f
c98 87 Vss 2.60675e-19
c99 81 Vss 0.00257188f
c100 76 Vss 7.28175e-19
c101 71 Vss 0.00117992f
c102 66 Vss 0.00174295f
c103 63 Vss 0.00812841f
c104 59 Vss 0.00683037f
c105 54 Vss 0.00816767f
c106 43 Vss 0.0342891f
c107 42 Vss 0.100071f
c108 33 Vss 0.0350852f
c109 32 Vss 0.0990713f
c110 14 Vss 0.00143493f
c111 11 Vss 0.378924f
c112 3 Vss 0.378636f
r113 142 146 0.349767
r114 141 142 5.50157
r115 137 146 0.306046
r116 130 144 0.494161
r117 129 141 0.652036
r118 125 144 0.128424
r119 123 133 0.652036
r120 123 124 10.1279
r121 119 143 0.0828784
r122 117 144 0.494161
r123 117 118 4.37625
r124 116 124 0.652036
r125 115 143 0.551426
r126 115 116 5.50157
r127 114 143 0.551426
r128 113 118 0.652036
r129 113 114 17.4633
r130 87 137 1.82344
r131 81 129 13.5872
r132 81 130 8.04396
r133 81 84 6.71025
r134 76 101 1.16709
r135 76 133 2.16729
r136 71 96 1.16709
r137 71 125 2.16729
r138 66 119 1.82344
r139 63 87 1.16709
r140 59 84 1.16709
r141 54 66 1.16709
r142 45 101 0.0476429
r143 43 45 1.45875
r144 42 46 0.652036
r145 42 45 1.45875
r146 39 43 0.652036
r147 35 96 0.0476429
r148 33 35 1.45875
r149 32 36 0.652036
r150 32 35 1.45875
r151 29 33 0.652036
r152 16 63 0.123773
r153 14 59 0.123773
r154 11 46 5.1348
r155 11 39 5.1348
r156 8 59 0.123773
r157 6 54 0.123773
r158 3 36 5.1348
r159 3 29 5.1348
.ends

.subckt PM_G4_XNOR2_N3_A 2 4 7 10 21 24 28 39 48 54 57 62 67 72 77 85 Vss
c54 85 Vss 5.19577e-19
c55 77 Vss 0.00107525f
c56 72 Vss 0.00526551f
c57 67 Vss 0.00394354f
c58 62 Vss 0.00276499f
c59 57 Vss 0.00595775f
c60 54 Vss 8.99321e-19
c61 48 Vss 0.126065f
c62 43 Vss 0.0296855f
c63 39 Vss 4.49964e-19
c64 28 Vss 0.152703f
c65 24 Vss 8.95828e-20
c66 21 Vss 0.173355f
c67 18 Vss 0.180502f
c68 16 Vss 0.0247918f
c69 10 Vss 0.176514f
c70 7 Vss 0.433917f
c71 4 Vss 0.193054f
r72 81 85 0.653045
r73 62 77 1.16709
r74 62 85 4.9014
r75 57 72 1.16709
r76 57 81 11.3366
r77 51 67 1.16709
r78 51 54 0.0364688
r79 47 72 0.0238214
r80 47 48 2.334
r81 44 47 2.20433
r82 39 77 0.404964
r83 33 48 0.00605528
r84 31 44 0.00605528
r85 29 43 0.494161
r86 28 30 0.652036
r87 28 29 4.84305
r88 25 43 0.128424
r89 24 67 0.0476429
r90 22 24 0.326018
r91 22 24 0.1167
r92 21 43 0.494161
r93 21 24 6.7686
r94 18 67 0.357321
r95 16 24 0.326018
r96 16 18 0.40845
r97 10 39 4.60965
r98 7 33 5.1348
r99 7 31 5.1348
r100 7 30 5.1348
r101 4 25 5.1348
r102 2 18 4.72635
.ends

.subckt PM_G4_XNOR2_N3_NET1 2 4 7 10 30 31 35 41 44 49 58 66 Vss
c34 66 Vss 2.27666e-19
c35 58 Vss 0.0070279f
c36 49 Vss 0.00633509f
c37 44 Vss 0.0011111f
c38 41 Vss 0.00508953f
c39 35 Vss 0.103132f
c40 31 Vss 0.128995f
c41 30 Vss 9.4155e-20
c42 10 Vss 0.290846f
c43 7 Vss 0.485246f
c44 4 Vss 0.00143493f
r45 62 66 0.653045
r46 49 58 1.16709
r47 49 66 12.9148
r48 44 62 3.37596
r49 41 44 1.16709
r50 33 35 1.70187
r51 30 58 0.0238214
r52 30 31 2.20433
r53 27 30 2.334
r54 25 35 0.17282
r55 24 31 0.00605528
r56 21 33 0.17282
r57 18 27 0.00605528
r58 10 21 8.34405
r59 7 25 7.002
r60 7 24 5.1348
r61 7 18 5.1348
r62 4 41 0.123773
r63 2 41 0.123773
.ends

.subckt PM_G4_XNOR2_N3_NET3 2 4 6 9 21 22 33 39 42 47 56 74 Vss
c47 74 Vss 3.98722e-19
c48 56 Vss 0.00391617f
c49 47 Vss 0.00744607f
c50 42 Vss 0.00230693f
c51 39 Vss 0.00508953f
c52 33 Vss 0.12548f
c53 22 Vss 0.0328697f
c54 21 Vss 0.175168f
c55 9 Vss 0.574903f
c56 6 Vss 0.200347f
c57 4 Vss 0.00143493f
r58 70 74 0.660011
r59 47 56 1.16709
r60 47 74 11.3611
r61 42 70 3.29261
r62 39 42 1.16709
r63 32 56 0.0238214
r64 32 33 2.26917
r65 29 32 2.26917
r66 26 33 0.00605528
r67 24 29 0.00605528
r68 21 23 0.652036
r69 21 22 4.84305
r70 18 22 0.652036
r71 9 26 5.1348
r72 9 24 5.1348
r73 9 23 10.0362
r74 6 18 5.54325
r75 4 39 0.123773
r76 2 39 0.123773
.ends

.subckt PM_G4_XNOR2_N3_B 2 4 7 10 19 20 28 31 33 37 38 48 52 55 58 61 Vss
c34 61 Vss 0.0283565f
c35 55 Vss 0.00145453f
c36 52 Vss 0.136463f
c37 48 Vss 0.0595773f
c38 38 Vss 0.0333783f
c39 37 Vss 0.0913542f
c40 33 Vss 0.0446983f
c41 31 Vss 8.50018e-20
c42 28 Vss 0.0899906f
c43 20 Vss 0.0348606f
c44 19 Vss 0.173355f
c45 10 Vss 0.264298f
c46 7 Vss 0.429172f
c47 4 Vss 0.180506f
c48 2 Vss 0.192541f
r49 55 61 1.16709
r50 55 58 0.0416786
r51 50 52 4.53833
r52 47 48 1.167
r53 42 52 0.00605528
r54 37 39 0.652036
r55 37 38 2.04225
r56 35 48 0.0685365
r57 34 50 0.00605528
r58 33 38 0.652036
r59 32 47 0.0685365
r60 32 33 1.69215
r61 31 61 0.181909
r62 29 61 0.494161
r63 29 31 0.1167
r64 28 47 0.5835
r65 28 31 3.55935
r66 23 61 0.128424
r67 23 61 0.40845
r68 22 61 0.181909
r69 20 22 6.7686
r70 19 61 0.494161
r71 19 22 0.1167
r72 16 20 0.652036
r73 10 39 7.5855
r74 7 42 5.1348
r75 7 35 5.1348
r76 7 34 5.1348
r77 4 61 4.72635
r78 2 16 5.1348
.ends

.subckt PM_G4_XNOR2_N3_Z 2 4 6 8 23 27 30 33 Vss
c28 30 Vss 0.0035978f
c29 27 Vss 0.00609752f
c30 23 Vss 0.00569635f
c31 8 Vss 0.00143493f
c32 6 Vss 0.00143493f
r33 33 35 5.29318
r34 30 33 6.66857
r35 27 35 1.16709
r36 23 30 1.16709
r37 8 27 0.123773
r38 6 23 0.123773
r39 4 27 0.123773
r40 2 23 0.123773
.ends

.subckt G4_XNOR2_N3  VDD VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI20.X0 N_NET1_XI20.X0_D N_VSS_XI20.X0_PGD N_B_XI20.X0_CG N_VSS_XI20.X0_PGD
+ N_VDD_XI20.X0_S TIGFET_HPNW12
XI24.X0 N_NET3_XI24.X0_D N_VDD_XI24.X0_PGD N_A_XI24.X0_CG N_VDD_XI24.X0_PGD
+ N_VSS_XI24.X0_S TIGFET_HPNW12
XI22.X0 N_NET1_XI22.X0_D N_VDD_XI22.X0_PGD N_B_XI22.X0_CG N_VDD_XI22.X0_PGD
+ N_VSS_XI22.X0_S TIGFET_HPNW12
XI26.X0 N_NET3_XI26.X0_D N_VSS_XI26.X0_PGD N_A_XI26.X0_CG N_VSS_XI26.X0_PGD
+ N_VDD_XI26.X0_S TIGFET_HPNW12
XI21.X0 N_Z_XI21.X0_D N_B_XI21.X0_PGD N_NET3_XI21.X0_CG N_B_XI21.X0_PGD
+ N_VSS_XI21.X0_S TIGFET_HPNW12
XI25.X0 N_Z_XI25.X0_D N_A_XI25.X0_PGD N_B_XI25.X0_CG N_A_XI25.X0_PGD
+ N_VDD_XI25.X0_S TIGFET_HPNW12
XI23.X0 N_Z_XI23.X0_D N_NET1_XI23.X0_PGD N_A_XI23.X0_CG N_NET1_XI23.X0_PGD
+ N_VSS_XI23.X0_S TIGFET_HPNW12
XI27.X0 N_Z_XI27.X0_D N_NET3_XI27.X0_PGD N_NET1_XI27.X0_CG N_NET3_XI27.X0_PGD
+ N_VDD_XI27.X0_S TIGFET_HPNW12
*
x_PM_G4_XNOR2_N3_VDD N_VDD_XI20.X0_S N_VDD_XI24.X0_PGD N_VDD_XI22.X0_PGD
+ N_VDD_XI26.X0_S N_VDD_XI25.X0_S N_VDD_XI27.X0_S N_VDD_c_9_p N_VDD_c_23_p
+ N_VDD_c_5_p N_VDD_c_89_p N_VDD_c_64_p N_VDD_c_11_p N_VDD_c_7_p N_VDD_c_12_p
+ N_VDD_c_6_p N_VDD_c_39_p N_VDD_c_13_p N_VDD_c_14_p N_VDD_c_43_p N_VDD_c_19_p
+ N_VDD_c_10_p N_VDD_c_17_p N_VDD_c_4_p N_VDD_c_53_p N_VDD_c_45_p N_VDD_c_59_p
+ N_VDD_c_36_p N_VDD_c_42_p VDD N_VDD_c_22_p N_VDD_c_18_p N_VDD_c_97_p Vss
+ PM_G4_XNOR2_N3_VDD
x_PM_G4_XNOR2_N3_VSS N_VSS_XI20.X0_PGD N_VSS_XI24.X0_S N_VSS_XI22.X0_S
+ N_VSS_XI26.X0_PGD N_VSS_XI21.X0_S N_VSS_XI23.X0_S N_VSS_c_107_n N_VSS_c_109_n
+ N_VSS_c_154_p N_VSS_c_111_n N_VSS_c_170_p N_VSS_c_113_n N_VSS_c_181_p
+ N_VSS_c_114_n N_VSS_c_117_n N_VSS_c_121_n N_VSS_c_125_n N_VSS_c_183_p
+ N_VSS_c_129_n N_VSS_c_133_n N_VSS_c_136_n N_VSS_c_139_n N_VSS_c_140_n
+ N_VSS_c_141_n N_VSS_c_142_n N_VSS_c_145_n N_VSS_c_146_n N_VSS_c_147_n
+ N_VSS_c_165_p N_VSS_c_148_n N_VSS_c_149_n VSS Vss PM_G4_XNOR2_N3_VSS
x_PM_G4_XNOR2_N3_A N_A_XI24.X0_CG N_A_XI26.X0_CG N_A_XI25.X0_PGD N_A_XI23.X0_CG
+ N_A_c_189_n N_A_c_191_n N_A_c_192_n N_A_c_215_p N_A_c_193_n A N_A_c_197_n
+ N_A_c_216_p N_A_c_200_n N_A_c_202_n N_A_c_214_p N_A_c_212_n Vss
+ PM_G4_XNOR2_N3_A
x_PM_G4_XNOR2_N3_NET1 N_NET1_XI20.X0_D N_NET1_XI22.X0_D N_NET1_XI23.X0_PGD
+ N_NET1_XI27.X0_CG N_NET1_c_263_n N_NET1_c_274_p N_NET1_c_267_p N_NET1_c_242_n
+ N_NET1_c_245_n N_NET1_c_249_n N_NET1_c_257_n N_NET1_c_258_n Vss
+ PM_G4_XNOR2_N3_NET1
x_PM_G4_XNOR2_N3_NET3 N_NET3_XI24.X0_D N_NET3_XI26.X0_D N_NET3_XI21.X0_CG
+ N_NET3_XI27.X0_PGD N_NET3_c_298_n N_NET3_c_314_p N_NET3_c_277_n N_NET3_c_278_n
+ N_NET3_c_279_n N_NET3_c_282_n N_NET3_c_285_n N_NET3_c_287_n Vss
+ PM_G4_XNOR2_N3_NET3
x_PM_G4_XNOR2_N3_B N_B_XI20.X0_CG N_B_XI22.X0_CG N_B_XI21.X0_PGD N_B_XI25.X0_CG
+ N_B_c_325_n N_B_c_338_n N_B_c_327_n N_B_c_328_n N_B_c_351_n N_B_c_347_n
+ N_B_c_340_n N_B_c_341_n N_B_c_329_n N_B_c_330_n B N_B_c_331_n Vss
+ PM_G4_XNOR2_N3_B
x_PM_G4_XNOR2_N3_Z N_Z_XI21.X0_D N_Z_XI25.X0_D N_Z_XI23.X0_D N_Z_XI27.X0_D
+ N_Z_c_367_n N_Z_c_357_n N_Z_c_362_n Z Vss PM_G4_XNOR2_N3_Z
cc_1 N_VDD_XI24.X0_PGD N_VSS_XI20.X0_PGD 2.9783e-19
cc_2 N_VDD_XI22.X0_PGD N_VSS_XI20.X0_PGD 0.0019598f
cc_3 N_VDD_XI24.X0_PGD N_VSS_XI26.X0_PGD 0.0019593f
cc_4 N_VDD_c_4_p N_VSS_XI26.X0_PGD 2.21956e-19
cc_5 N_VDD_c_5_p N_VSS_c_107_n 0.0019598f
cc_6 N_VDD_c_6_p N_VSS_c_107_n 3.89167e-19
cc_7 N_VDD_c_7_p N_VSS_c_109_n 3.80615e-19
cc_8 N_VDD_c_6_p N_VSS_c_109_n 3.89167e-19
cc_9 N_VDD_c_9_p N_VSS_c_111_n 0.0019593f
cc_10 N_VDD_c_10_p N_VSS_c_111_n 3.89167e-19
cc_11 N_VDD_c_11_p N_VSS_c_113_n 3.47417e-19
cc_12 N_VDD_c_12_p N_VSS_c_114_n 0.00187494f
cc_13 N_VDD_c_13_p N_VSS_c_114_n 4.32036e-19
cc_14 N_VDD_c_14_p N_VSS_c_114_n 3.5277e-19
cc_15 N_VDD_c_7_p N_VSS_c_117_n 4.35319e-19
cc_16 N_VDD_c_6_p N_VSS_c_117_n 0.00161703f
cc_17 N_VDD_c_17_p N_VSS_c_117_n 8.66259e-19
cc_18 N_VDD_c_18_p N_VSS_c_117_n 3.48267e-19
cc_19 N_VDD_c_19_p N_VSS_c_121_n 9.53113e-19
cc_20 N_VDD_c_10_p N_VSS_c_121_n 0.00161703f
cc_21 N_VDD_c_4_p N_VSS_c_121_n 0.00227183f
cc_22 N_VDD_c_22_p N_VSS_c_121_n 3.48267e-19
cc_23 N_VDD_c_23_p N_VSS_c_125_n 2.36481e-19
cc_24 N_VDD_c_6_p N_VSS_c_125_n 0.00538298f
cc_25 N_VDD_c_4_p N_VSS_c_125_n 2.5578e-19
cc_26 N_VDD_c_18_p N_VSS_c_125_n 9.58524e-19
cc_27 N_VDD_c_7_p N_VSS_c_129_n 3.66936e-19
cc_28 N_VDD_c_6_p N_VSS_c_129_n 2.26455e-19
cc_29 N_VDD_c_17_p N_VSS_c_129_n 3.99794e-19
cc_30 N_VDD_c_18_p N_VSS_c_129_n 6.489e-19
cc_31 N_VDD_c_10_p N_VSS_c_133_n 2.26455e-19
cc_32 N_VDD_c_4_p N_VSS_c_133_n 9.55322e-19
cc_33 N_VDD_c_22_p N_VSS_c_133_n 6.46219e-19
cc_34 N_VDD_c_7_p N_VSS_c_136_n 0.00378845f
cc_35 N_VDD_c_12_p N_VSS_c_136_n 0.00917884f
cc_36 N_VDD_c_36_p N_VSS_c_136_n 0.0010706f
cc_37 N_VDD_c_12_p N_VSS_c_139_n 0.00404533f
cc_38 N_VDD_c_6_p N_VSS_c_140_n 0.00348469f
cc_39 N_VDD_c_39_p N_VSS_c_141_n 0.00107963f
cc_40 N_VDD_c_14_p N_VSS_c_142_n 0.00356332f
cc_41 N_VDD_c_10_p N_VSS_c_142_n 0.00615517f
cc_42 N_VDD_c_42_p N_VSS_c_142_n 9.37919e-19
cc_43 N_VDD_c_43_p N_VSS_c_145_n 0.00106367f
cc_44 N_VDD_c_6_p N_VSS_c_146_n 0.00468936f
cc_45 N_VDD_c_45_p N_VSS_c_147_n 9.00324e-19
cc_46 N_VDD_c_12_p N_VSS_c_148_n 9.16632e-19
cc_47 N_VDD_c_6_p N_VSS_c_149_n 7.74609e-19
cc_48 N_VDD_c_4_p N_A_XI25.X0_PGD 2.05446e-19
cc_49 N_VDD_XI24.X0_PGD N_A_c_189_n 4.09718e-19
cc_50 N_VDD_XI22.X0_PGD N_A_c_189_n 2.22577e-19
cc_51 N_VDD_c_22_p N_A_c_191_n 5.33384e-19
cc_52 N_VDD_XI22.X0_PGD N_A_c_192_n 2.22577e-19
cc_53 N_VDD_c_53_p N_A_c_193_n 6.08999e-19
cc_54 N_VDD_c_12_p A 5.04211e-19
cc_55 N_VDD_c_19_p A 2.95248e-19
cc_56 N_VDD_c_22_p A 2.15082e-19
cc_57 N_VDD_c_4_p N_A_c_197_n 0.00289813f
cc_58 N_VDD_c_53_p N_A_c_197_n 0.00191817f
cc_59 N_VDD_c_59_p N_A_c_197_n 3.22661e-19
cc_60 N_VDD_c_12_p N_A_c_200_n 6.25289e-19
cc_61 N_VDD_c_19_p N_A_c_200_n 2.28697e-19
cc_62 N_VDD_c_4_p N_A_c_202_n 9.84209e-19
cc_63 N_VDD_c_53_p N_A_c_202_n 2.68554e-19
cc_64 N_VDD_c_64_p N_NET1_c_242_n 3.43419e-19
cc_65 N_VDD_c_6_p N_NET1_c_242_n 2.74986e-19
cc_66 N_VDD_c_13_p N_NET1_c_242_n 3.72199e-19
cc_67 N_VDD_c_64_p N_NET1_c_245_n 3.48267e-19
cc_68 N_VDD_c_7_p N_NET1_c_245_n 2.34601e-19
cc_69 N_VDD_c_6_p N_NET1_c_245_n 2.9533e-19
cc_70 N_VDD_c_13_p N_NET1_c_245_n 5.226e-19
cc_71 N_VDD_c_17_p N_NET1_c_249_n 0.00122163f
cc_72 N_VDD_c_59_p N_NET3_XI27.X0_PGD 4.14305e-19
cc_73 N_VDD_c_53_p N_NET3_c_277_n 8.42825e-19
cc_74 N_VDD_c_11_p N_NET3_c_278_n 3.43419e-19
cc_75 N_VDD_c_11_p N_NET3_c_279_n 3.48267e-19
cc_76 N_VDD_c_10_p N_NET3_c_279_n 3.21336e-19
cc_77 N_VDD_c_4_p N_NET3_c_279_n 0.00123864f
cc_78 N_VDD_c_4_p N_NET3_c_282_n 0.00123016f
cc_79 N_VDD_c_53_p N_NET3_c_282_n 0.00291325f
cc_80 N_VDD_c_59_p N_NET3_c_282_n 7.77543e-19
cc_81 N_VDD_c_53_p N_NET3_c_285_n 0.00118178f
cc_82 N_VDD_c_59_p N_NET3_c_285_n 3.66936e-19
cc_83 N_VDD_c_19_p N_NET3_c_287_n 3.02266e-19
cc_84 N_VDD_c_12_p N_B_XI20.X0_CG 3.50093e-19
cc_85 N_VDD_XI22.X0_PGD N_B_XI21.X0_PGD 0.00190378f
cc_86 N_VDD_XI24.X0_PGD N_B_c_325_n 2.22577e-19
cc_87 N_VDD_XI22.X0_PGD N_B_c_325_n 4.09718e-19
cc_88 N_VDD_XI22.X0_PGD N_B_c_327_n 4.09718e-19
cc_89 N_VDD_c_89_p N_B_c_328_n 5.7019e-19
cc_90 N_VDD_c_23_p N_B_c_329_n 0.00168656f
cc_91 N_VDD_c_18_p N_B_c_330_n 2.15082e-19
cc_92 N_VDD_c_17_p N_B_c_331_n 2.26584e-19
cc_93 N_VDD_c_11_p N_Z_c_357_n 3.43419e-19
cc_94 N_VDD_c_4_p N_Z_c_357_n 3.48267e-19
cc_95 N_VDD_c_53_p N_Z_c_357_n 2.74986e-19
cc_96 N_VDD_c_45_p N_Z_c_357_n 3.72199e-19
cc_97 N_VDD_c_97_p N_Z_c_357_n 3.43419e-19
cc_98 N_VDD_c_11_p N_Z_c_362_n 3.48267e-19
cc_99 N_VDD_c_4_p N_Z_c_362_n 4.85404e-19
cc_100 N_VDD_c_53_p N_Z_c_362_n 4.9751e-19
cc_101 N_VDD_c_45_p N_Z_c_362_n 8.21216e-19
cc_102 N_VDD_c_97_p N_Z_c_362_n 3.48267e-19
cc_103 N_VSS_XI26.X0_PGD N_A_XI25.X0_PGD 0.00164979f
cc_104 N_VSS_XI20.X0_PGD N_A_c_189_n 2.22577e-19
cc_105 N_VSS_XI26.X0_PGD N_A_c_189_n 4.09718e-19
cc_106 N_VSS_XI26.X0_PGD N_A_c_192_n 4.09718e-19
cc_107 N_VSS_c_154_p N_A_c_193_n 0.00164979f
cc_108 N_VSS_c_121_n N_A_c_197_n 3.87149e-19
cc_109 N_VSS_c_136_n N_A_c_197_n 6.21456e-19
cc_110 N_VSS_c_133_n N_A_c_202_n 6.52904e-19
cc_111 N_VSS_c_146_n N_A_c_212_n 5.04853e-19
cc_112 N_VSS_c_113_n N_NET1_c_242_n 3.43419e-19
cc_113 N_VSS_c_125_n N_NET1_c_242_n 3.48267e-19
cc_114 N_VSS_c_113_n N_NET1_c_245_n 3.48267e-19
cc_115 N_VSS_c_125_n N_NET1_c_245_n 0.00164479f
cc_116 N_VSS_c_125_n N_NET1_c_249_n 0.00162978f
cc_117 N_VSS_c_146_n N_NET1_c_249_n 0.0181004f
cc_118 N_VSS_c_165_p N_NET1_c_249_n 0.00121213f
cc_119 N_VSS_c_125_n N_NET1_c_257_n 2.78343e-19
cc_120 N_VSS_c_117_n N_NET1_c_258_n 0.00198862f
cc_121 N_VSS_c_136_n N_NET1_c_258_n 0.00136675f
cc_122 N_VSS_c_146_n N_NET1_c_258_n 0.00168829f
cc_123 N_VSS_c_170_p N_NET3_c_278_n 3.43419e-19
cc_124 N_VSS_c_170_p N_NET3_c_279_n 3.48267e-19
cc_125 N_VSS_c_114_n N_NET3_c_279_n 0.0011211f
cc_126 N_VSS_c_139_n N_NET3_c_279_n 6.33709e-19
cc_127 N_VSS_c_121_n N_NET3_c_282_n 0.00131985f
cc_128 N_VSS_c_142_n N_NET3_c_287_n 4.84133e-19
cc_129 N_VSS_XI20.X0_PGD N_B_c_325_n 4.09718e-19
cc_130 N_VSS_XI26.X0_PGD N_B_c_325_n 2.22577e-19
cc_131 N_VSS_XI26.X0_PGD N_B_c_327_n 2.22577e-19
cc_132 N_VSS_c_125_n N_B_c_329_n 2.44335e-19
cc_133 N_VSS_c_113_n N_Z_c_367_n 3.43419e-19
cc_134 N_VSS_c_181_p N_Z_c_367_n 3.43419e-19
cc_135 N_VSS_c_125_n N_Z_c_367_n 3.48267e-19
cc_136 N_VSS_c_183_p N_Z_c_367_n 3.48267e-19
cc_137 N_VSS_c_113_n N_Z_c_362_n 3.48267e-19
cc_138 N_VSS_c_181_p N_Z_c_362_n 3.48267e-19
cc_139 N_VSS_c_125_n N_Z_c_362_n 8.69457e-19
cc_140 N_VSS_c_183_p N_Z_c_362_n 5.71987e-19
cc_141 N_A_XI23.X0_CG N_NET1_XI23.X0_PGD 5.00154e-19
cc_142 N_A_c_214_p N_NET1_XI23.X0_PGD 0.0013363f
cc_143 N_A_c_215_p N_NET1_c_263_n 5.8445e-19
cc_144 N_A_c_216_p N_NET1_c_249_n 0.0020999f
cc_145 N_A_c_212_n N_NET1_c_249_n 6.74055e-19
cc_146 N_A_c_214_p N_NET3_XI21.X0_CG 2.18475e-19
cc_147 N_A_XI25.X0_PGD N_NET3_XI27.X0_PGD 0.00173934f
cc_148 N_A_c_192_n N_NET3_XI27.X0_PGD 3.14428e-19
cc_149 N_A_c_214_p N_NET3_XI27.X0_PGD 4.34237e-19
cc_150 N_A_XI25.X0_PGD N_NET3_c_298_n 4.64512e-19
cc_151 N_A_c_193_n N_NET3_c_277_n 0.00173934f
cc_152 N_A_c_189_n N_NET3_c_278_n 6.35441e-19
cc_153 N_A_c_197_n N_NET3_c_279_n 0.00122226f
cc_154 N_A_c_197_n N_NET3_c_282_n 0.00256249f
cc_155 N_A_c_216_p N_NET3_c_282_n 0.00124966f
cc_156 N_A_c_202_n N_NET3_c_282_n 3.44698e-19
cc_157 N_A_c_197_n N_NET3_c_285_n 3.44698e-19
cc_158 N_A_c_202_n N_NET3_c_285_n 6.70706e-19
cc_159 N_A_c_192_n N_B_XI25.X0_CG 0.003858f
cc_160 N_A_c_189_n N_B_c_325_n 0.00503082f
cc_161 N_A_c_200_n N_B_c_338_n 7.5077e-19
cc_162 N_A_c_192_n N_B_c_327_n 0.00270268f
cc_163 N_A_c_192_n N_B_c_340_n 0.00358164f
cc_164 N_A_c_192_n N_B_c_341_n 2.04018e-19
cc_165 N_A_c_212_n N_B_c_330_n 2.24721e-19
cc_166 N_A_c_189_n N_B_c_331_n 8.36919e-19
cc_167 N_A_c_197_n N_Z_c_362_n 0.00453915f
cc_168 N_A_c_216_p N_Z_c_362_n 0.00285282f
cc_169 N_A_c_214_p N_Z_c_362_n 9.79999e-19
cc_170 N_NET1_XI23.X0_PGD N_NET3_XI21.X0_CG 3.25363e-19
cc_171 N_NET1_c_267_p N_NET3_XI27.X0_PGD 0.00866857f
cc_172 N_NET1_XI23.X0_PGD N_NET3_c_298_n 0.00335065f
cc_173 N_NET1_c_242_n N_NET3_c_278_n 2.56771e-19
cc_174 N_NET1_XI23.X0_PGD N_B_XI21.X0_PGD 0.00216073f
cc_175 N_NET1_XI27.X0_CG N_B_XI25.X0_CG 2.72501e-19
cc_176 N_NET1_c_242_n N_B_c_325_n 6.35441e-19
cc_177 N_NET1_c_267_p N_B_c_347_n 2.72501e-19
cc_178 N_NET1_c_274_p N_B_c_329_n 0.00193498f
cc_179 N_NET1_c_249_n N_Z_c_362_n 3.17674e-19
cc_180 N_NET3_XI21.X0_CG N_B_XI21.X0_PGD 0.00200964f
cc_181 N_NET3_c_298_n N_B_XI21.X0_PGD 0.00163867f
cc_182 N_NET3_XI27.X0_PGD N_B_c_351_n 3.23792e-19
cc_183 N_NET3_c_314_p N_B_c_351_n 5.75226e-19
cc_184 N_NET3_XI27.X0_PGD N_B_c_347_n 0.00310335f
cc_185 N_NET3_c_314_p N_B_c_347_n 0.00201276f
cc_186 N_NET3_c_314_p N_B_c_341_n 0.00200964f
cc_187 N_NET3_c_298_n N_Z_c_367_n 6.58359e-19
cc_188 N_NET3_c_298_n N_Z_c_357_n 2.51847e-19
cc_189 N_NET3_XI27.X0_PGD N_Z_c_362_n 0.00129454f
cc_190 N_NET3_c_298_n N_Z_c_362_n 2.39178e-19
cc_191 N_NET3_c_282_n N_Z_c_362_n 2.33494e-19
cc_192 N_B_c_347_n N_Z_c_362_n 9.47639e-19
*
.ends
*
*
.subckt XNOR2_HPNW12 A B Y VDD VSS
xgate (VDD VSS A B Y) G4_XNOR2_N3
.ends
*
* File: G5_XNOR3_N3.pex.netlist
* Created: Mon Mar 28 16:13:50 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XNOR3_N3_VDD 2 5 9 12 14 17 34 35 44 45 54 55 65 69 74 77 79 80 81
+ 84 86 87 90 93 96 98 102 104 108 112 114 116 117 119 125 134 139 Vss
c113 139 Vss 0.0048986f
c114 134 Vss 0.00495479f
c115 125 Vss 0.00563771f
c116 117 Vss 2.39889e-19
c117 116 Vss 4.92173e-19
c118 115 Vss 5.21614e-19
c119 114 Vss 4.52364e-19
c120 112 Vss 0.0017155f
c121 110 Vss 0.00173699f
c122 108 Vss 6.49327e-19
c123 104 Vss 0.00471178f
c124 102 Vss 0.0010418f
c125 98 Vss 0.00587581f
c126 96 Vss 0.00147489f
c127 93 Vss 0.00334883f
c128 90 Vss 0.00547221f
c129 87 Vss 8.67855e-19
c130 86 Vss 0.00654417f
c131 84 Vss 0.00154142f
c132 81 Vss 8.68392e-19
c133 80 Vss 0.00938293f
c134 79 Vss 0.0116507f
c135 77 Vss 0.00304889f
c136 74 Vss 0.00785043f
c137 69 Vss 0.00836757f
c138 65 Vss 0.00811483f
c139 55 Vss 0.0356247f
c140 54 Vss 0.10084f
c141 45 Vss 0.0356281f
c142 44 Vss 0.101312f
c143 35 Vss 0.0346562f
c144 34 Vss 0.0991017f
c145 17 Vss 0.378772f
c146 9 Vss 0.379175f
c147 5 Vss 0.383323f
r148 110 119 0.326018
r149 110 112 6.16843
r150 108 139 1.16709
r151 106 108 2.16729
r152 105 117 0.494161
r153 104 119 0.326018
r154 104 105 7.46046
r155 102 134 1.16709
r156 100 117 0.128424
r157 100 102 2.16729
r158 99 116 0.494161
r159 98 106 0.652036
r160 98 99 10.3363
r161 94 115 0.0828784
r162 94 96 2.00578
r163 93 116 0.128424
r164 92 115 0.551426
r165 92 93 5.50157
r166 90 125 1.16709
r167 88 115 0.551426
r168 88 90 7.66886
r169 86 116 0.494161
r170 86 87 10.1279
r171 82 114 0.0828784
r172 82 84 1.82344
r173 80 117 0.494161
r174 80 81 15.8795
r175 79 87 0.652036
r176 78 114 0.551426
r177 78 79 18.3386
r178 77 114 0.551426
r179 76 81 0.652036
r180 76 77 5.50157
r181 74 112 1.16709
r182 69 96 1.16709
r183 65 84 1.16709
r184 57 139 0.0476429
r185 55 57 1.45875
r186 54 58 0.652036
r187 54 57 1.45875
r188 51 55 0.652036
r189 47 134 0.0476429
r190 45 47 1.45875
r191 44 48 0.652036
r192 44 47 1.45875
r193 41 45 0.652036
r194 37 125 0.238214
r195 35 37 1.45875
r196 34 38 0.652036
r197 34 37 1.45875
r198 31 35 0.652036
r199 17 58 5.1348
r200 17 51 5.1348
r201 14 74 0.123773
r202 12 69 0.123773
r203 9 48 5.1348
r204 9 41 5.1348
r205 5 38 5.1348
r206 5 31 5.1348
r207 2 65 0.123773
.ends

.subckt PM_G5_XNOR3_N3_C 2 4 6 8 17 20 23 32 37 40 44 47 52 57 84 92 98 Vss
c49 98 Vss 3.10785e-19
c50 92 Vss 0.00560641f
c51 84 Vss 0.00950787f
c52 57 Vss 0.004971f
c53 52 Vss 7.31067e-19
c54 47 Vss 0.00104925f
c55 40 Vss 0.00163759f
c56 37 Vss 0.0082356f
c57 32 Vss 0.00958317f
c58 23 Vss 2.04877e-19
c59 20 Vss 0.221837f
c60 17 Vss 0.180502f
c61 15 Vss 0.0247918f
c62 4 Vss 0.188411f
r63 93 98 0.441572
r64 92 94 0.655813
r65 92 93 9.04425
r66 88 98 0.174814
r67 84 98 0.441572
r68 52 94 3.33429
r69 47 88 3.33429
r70 40 57 1.16709
r71 40 84 22.1365
r72 40 44 0.0833571
r73 37 52 1.16709
r74 32 47 1.16709
r75 23 57 0.0476429
r76 21 23 0.326018
r77 21 23 0.1167
r78 20 24 0.652036
r79 20 23 6.7686
r80 17 57 0.357321
r81 15 23 0.326018
r82 15 17 0.40845
r83 8 37 0.123773
r84 6 32 0.123773
r85 4 24 5.1348
r86 2 17 4.72635
.ends

.subckt PM_G5_XNOR3_N3_VSS 3 6 8 11 15 18 34 37 44 45 54 55 57 66 70 73 78 83 88
+ 93 96 99 108 113 122 124 125 126 131 132 137 149 153 154 155 Vss
c122 155 Vss 3.75522e-19
c123 154 Vss 3.91906e-19
c124 153 Vss 4.4306e-19
c125 149 Vss 3.17876e-19
c126 137 Vss 0.00359616f
c127 132 Vss 8.45126e-19
c128 131 Vss 0.00635332f
c129 126 Vss 8.42189e-19
c130 125 Vss 0.0059194f
c131 124 Vss 0.00452138f
c132 122 Vss 0.00375531f
c133 113 Vss 0.00410359f
c134 108 Vss 0.00419612f
c135 99 Vss 0.00605485f
c136 96 Vss 0.00346991f
c137 93 Vss 0.00310291f
c138 88 Vss 2.34373e-19
c139 83 Vss 0.00134516f
c140 78 Vss 0.0023966f
c141 73 Vss 0.00367309f
c142 70 Vss 0.0100681f
c143 66 Vss 0.00715185f
c144 57 Vss 9.33833e-20
c145 55 Vss 0.0347733f
c146 54 Vss 0.0999406f
c147 45 Vss 0.035088f
c148 44 Vss 0.0994129f
c149 37 Vss 5.39995e-20
c150 35 Vss 0.0349058f
c151 34 Vss 0.100344f
c152 15 Vss 0.379275f
c153 11 Vss 0.379887f
c154 8 Vss 0.00143493f
c155 3 Vss 0.3841f
r156 147 149 0.416786
r157 143 155 0.494161
r158 139 155 0.128424
r159 138 154 0.494161
r160 137 147 0.652036
r161 137 138 7.46046
r162 133 154 0.128424
r163 131 155 0.494161
r164 131 132 15.8795
r165 127 153 0.0828784
r166 125 154 0.494161
r167 125 126 13.0037
r168 124 132 0.652036
r169 123 153 0.551426
r170 123 124 13.8373
r171 122 153 0.551426
r172 121 126 0.652036
r173 121 122 10.0029
r174 96 143 8.04396
r175 93 96 6.75193
r176 88 113 1.16709
r177 88 149 1.7505
r178 83 108 1.16709
r179 83 139 2.16729
r180 78 133 6.16843
r181 73 99 1.16709
r182 73 127 4.33978
r183 70 93 1.16709
r184 66 78 1.16709
r185 57 113 0.0476429
r186 55 57 1.45875
r187 54 58 0.652036
r188 54 57 1.45875
r189 51 55 0.652036
r190 47 108 0.0476429
r191 45 47 1.45875
r192 44 48 0.652036
r193 44 47 1.45875
r194 41 45 0.652036
r195 37 99 0.238214
r196 35 37 1.45875
r197 34 38 0.652036
r198 34 37 1.45875
r199 31 35 0.652036
r200 18 70 0.123773
r201 15 58 5.1348
r202 15 51 5.1348
r203 11 48 5.1348
r204 11 41 5.1348
r205 8 66 0.123773
r206 6 66 0.123773
r207 3 38 5.1348
r208 3 31 5.1348
.ends

.subckt PM_G5_XNOR3_N3_CI 2 4 6 8 23 26 31 34 39 44 79 80 85 91 Vss
c47 91 Vss 2.55674e-19
c48 85 Vss 0.00650738f
c49 80 Vss 3.61784e-19
c50 79 Vss 0.00547357f
c51 44 Vss 7.31067e-19
c52 39 Vss 7.72278e-19
c53 34 Vss 0.00616608f
c54 31 Vss 0.00967911f
c55 26 Vss 0.00811165f
c56 23 Vss 0.00522928f
c57 4 Vss 0.00143493f
r58 86 91 0.441572
r59 85 87 0.655813
r60 85 86 9.04425
r61 81 91 0.174814
r62 79 91 0.441572
r63 79 80 19.1096
r64 75 80 0.655813
r65 44 87 3.33429
r66 39 81 3.33429
r67 34 75 16.1713
r68 31 44 1.16709
r69 26 39 1.16709
r70 23 34 1.16709
r71 8 31 0.123773
r72 6 26 0.123773
r73 4 23 0.123773
r74 2 23 0.123773
.ends

.subckt PM_G5_XNOR3_N3_A 2 4 7 11 24 44 45 49 51 54 56 57 60 65 66 69 74 Vss
c69 74 Vss 0.00565895f
c70 69 Vss 0.00509443f
c71 66 Vss 0.00618081f
c72 65 Vss 7.10913e-19
c73 57 Vss 8.70991e-19
c74 56 Vss 6.16621e-19
c75 54 Vss 0.00573533f
c76 51 Vss 0.00643922f
c77 49 Vss 0.135088f
c78 45 Vss 0.127808f
c79 44 Vss 1.14131e-19
c80 24 Vss 0.217341f
c81 21 Vss 0.18375f
c82 19 Vss 0.0247918f
c83 7 Vss 1.43795f
c84 4 Vss 0.194116f
r85 65 74 1.16709
r86 65 66 0.531835
r87 62 69 1.16709
r88 60 62 0.125036
r89 57 60 0.708536
r90 56 66 10.4613
r91 53 56 0.652036
r92 53 54 10.503
r93 52 57 0.0685365
r94 51 54 0.652036
r95 51 52 10.2113
r96 47 49 4.53833
r97 44 74 0.0238214
r98 44 45 2.26917
r99 41 44 2.26917
r100 36 49 0.00605528
r101 35 45 0.00605528
r102 32 47 0.00605528
r103 31 41 0.00605528
r104 27 69 0.0952857
r105 25 27 0.326018
r106 25 27 0.1167
r107 24 28 0.652036
r108 24 27 6.7686
r109 21 27 0.3335
r110 19 27 0.326018
r111 19 21 0.2334
r112 11 36 5.1348
r113 11 32 5.1348
r114 7 11 17.9718
r115 7 35 5.1348
r116 7 11 17.9718
r117 7 31 5.1348
r118 4 28 5.1348
r119 2 21 4.9014
.ends

.subckt PM_G5_XNOR3_N3_BI 2 4 6 8 16 23 29 32 37 42 51 56 64 65 68 77 82 83 Vss
c67 83 Vss 7.14146e-20
c68 82 Vss 6.9543e-19
c69 77 Vss 9.4202e-19
c70 68 Vss 6.59929e-19
c71 65 Vss 3.58032e-19
c72 64 Vss 0.00251452f
c73 56 Vss 0.00269072f
c74 51 Vss 0.0023082f
c75 42 Vss 0.00171238f
c76 37 Vss 4.65964e-19
c77 32 Vss 0.00208283f
c78 29 Vss 0.00520899f
c79 23 Vss 9.01088e-20
c80 16 Vss 0.166484f
c81 8 Vss 0.166484f
c82 4 Vss 0.00143493f
r83 81 83 0.65409
r84 81 82 3.42052
r85 77 82 0.652979
r86 68 77 2.03284
r87 66 68 2.00057
r88 64 66 0.652036
r89 64 65 13.2121
r90 60 65 0.652036
r91 42 56 1.16709
r92 42 83 2.00578
r93 37 51 1.16709
r94 37 68 0.0416786
r95 32 60 5.62661
r96 29 32 1.16709
r97 23 56 0.50025
r98 16 51 0.50025
r99 8 23 4.37625
r100 6 16 4.37625
r101 4 29 0.123773
r102 2 29 0.123773
.ends

.subckt PM_G5_XNOR3_N3_AI 2 4 7 11 31 37 43 46 51 60 68 Vss
c46 68 Vss 2.68274e-19
c47 60 Vss 0.00659076f
c48 51 Vss 0.00468816f
c49 46 Vss 8.13811e-19
c50 43 Vss 0.00461167f
c51 37 Vss 0.12791f
c52 31 Vss 0.134438f
c53 7 Vss 1.42501f
c54 4 Vss 0.00143493f
r55 64 68 0.655813
r56 51 60 1.16709
r57 51 68 12.0347
r58 46 64 3.33429
r59 43 46 1.16709
r60 36 60 0.0238214
r61 36 37 2.334
r62 33 36 2.20433
r63 29 31 4.53833
r64 26 37 0.00605528
r65 25 31 0.00605528
r66 22 33 0.00605528
r67 21 29 0.00605528
r68 11 26 5.1348
r69 11 22 5.1348
r70 7 11 17.9718
r71 7 25 5.1348
r72 7 11 17.9718
r73 7 21 5.1348
r74 4 43 0.123773
r75 2 43 0.123773
.ends

.subckt PM_G5_XNOR3_N3_B 2 4 6 8 16 17 24 31 41 44 49 54 59 65 69 76 77 Vss
c63 77 Vss 3.11913e-19
c64 76 Vss 9.9238e-19
c65 69 Vss 0.00389578f
c66 65 Vss 0.00255458f
c67 59 Vss 0.00150469f
c68 54 Vss 0.00172736f
c69 49 Vss 0.00131253f
c70 44 Vss 1.53364e-19
c71 41 Vss 3.86756e-19
c72 31 Vss 0.166484f
c73 24 Vss 8.82658e-20
c74 20 Vss 0.0247918f
c75 17 Vss 0.0339179f
c76 16 Vss 0.186033f
c77 6 Vss 0.166669f
c78 4 Vss 0.177261f
c79 2 Vss 0.191454f
r80 76 77 0.655813
r81 75 76 4.04282
r82 69 75 0.653045
r83 59 62 0.35
r84 49 65 1.16709
r85 49 77 2.00578
r86 44 59 1.16709
r87 44 69 2.1395
r88 41 54 1.16709
r89 41 44 10.7364
r90 36 54 0.309679
r91 31 65 0.50025
r92 28 62 0.452607
r93 24 54 0.214393
r94 20 36 0.326018
r95 20 24 0.75855
r96 17 36 6.7686
r97 16 36 0.326018
r98 16 36 0.1167
r99 13 17 0.652036
r100 8 31 4.37625
r101 6 28 4.2012
r102 4 24 4.37625
r103 2 13 5.1348
.ends

.subckt PM_G5_XNOR3_N3_Z 2 4 6 8 23 27 30 33 Vss
c30 30 Vss 0.00380939f
c31 27 Vss 0.00807893f
c32 23 Vss 0.00720799f
c33 8 Vss 0.00143493f
c34 6 Vss 0.00143493f
r35 33 35 6.33514
r36 30 33 6.50186
r37 27 35 1.16709
r38 23 30 1.16709
r39 8 27 0.123773
r40 6 23 0.123773
r41 4 27 0.123773
r42 2 23 0.123773
.ends

.subckt G5_XNOR3_N3  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI22.X0 N_CI_XI22.X0_D N_VSS_XI22.X0_PGD N_C_XI22.X0_CG N_VSS_XI22.X0_PGD
+ N_VDD_XI22.X0_S TIGFET_HPNW12
XI26.X0 N_CI_XI26.X0_D N_VDD_XI26.X0_PGD N_C_XI26.X0_CG N_VDD_XI26.X0_PGD
+ N_VSS_XI26.X0_S TIGFET_HPNW12
XI25.X0 N_BI_XI25.X0_D N_VDD_XI25.X0_PGD N_B_XI25.X0_CG N_VDD_XI25.X0_PGD
+ N_VSS_XI25.X0_S TIGFET_HPNW12
XI21.X0 N_AI_XI21.X0_D N_VSS_XI21.X0_PGD N_A_XI21.X0_CG N_VSS_XI21.X0_PGD
+ N_VDD_XI21.X0_S TIGFET_HPNW12
XI23.X0 N_BI_XI23.X0_D N_VSS_XI23.X0_PGD N_B_XI23.X0_CG N_VSS_XI23.X0_PGD
+ N_VDD_XI23.X0_S TIGFET_HPNW12
XI24.X0 N_AI_XI24.X0_D N_VDD_XI24.X0_PGD N_A_XI24.X0_CG N_VDD_XI24.X0_PGD
+ N_VSS_XI24.X0_S TIGFET_HPNW12
XI31.X0 N_Z_XI31.X0_D N_AI_XI31.X0_PGD N_B_XI31.X0_CG N_AI_XI31.X0_PGD
+ N_C_XI31.X0_S TIGFET_HPNW12
XI27.X0 N_Z_XI27.X0_D N_AI_XI27.X0_PGD N_BI_XI27.X0_CG N_AI_XI27.X0_PGD
+ N_CI_XI27.X0_S TIGFET_HPNW12
XI29.X0 N_Z_XI29.X0_D N_A_XI29.X0_PGD N_BI_XI29.X0_CG N_A_XI29.X0_PGD
+ N_C_XI29.X0_S TIGFET_HPNW12
XI28.X0 N_Z_XI28.X0_D N_A_XI28.X0_PGD N_B_XI28.X0_CG N_A_XI28.X0_PGD
+ N_CI_XI28.X0_S TIGFET_HPNW12
*
x_PM_G5_XNOR3_N3_VDD N_VDD_XI22.X0_S N_VDD_XI26.X0_PGD N_VDD_XI25.X0_PGD
+ N_VDD_XI21.X0_S N_VDD_XI23.X0_S N_VDD_XI24.X0_PGD N_VDD_c_112_p N_VDD_c_19_p
+ N_VDD_c_24_p N_VDD_c_4_p N_VDD_c_102_p N_VDD_c_20_p N_VDD_c_78_p N_VDD_c_103_p
+ N_VDD_c_6_p N_VDD_c_7_p N_VDD_c_13_p N_VDD_c_5_p N_VDD_c_64_p N_VDD_c_29_p
+ N_VDD_c_65_p N_VDD_c_69_p N_VDD_c_30_p N_VDD_c_16_p N_VDD_c_66_p N_VDD_c_21_p
+ N_VDD_c_10_p N_VDD_c_25_p N_VDD_c_37_p N_VDD_c_11_p N_VDD_c_60_p N_VDD_c_68_p
+ N_VDD_c_72_p VDD N_VDD_c_2_p N_VDD_c_42_p N_VDD_c_38_p Vss PM_G5_XNOR3_N3_VDD
x_PM_G5_XNOR3_N3_C N_C_XI22.X0_CG N_C_XI26.X0_CG N_C_XI31.X0_S N_C_XI29.X0_S
+ N_C_c_129_p N_C_c_116_n N_C_c_126_p N_C_c_119_n N_C_c_157_p N_C_c_120_n C
+ N_C_c_127_p N_C_c_159_p N_C_c_122_n N_C_c_123_n N_C_c_143_p N_C_c_148_p Vss
+ PM_G5_XNOR3_N3_C
x_PM_G5_XNOR3_N3_VSS N_VSS_XI22.X0_PGD N_VSS_XI26.X0_S N_VSS_XI25.X0_S
+ N_VSS_XI21.X0_PGD N_VSS_XI23.X0_PGD N_VSS_XI24.X0_S N_VSS_c_170_n
+ N_VSS_c_230_n N_VSS_c_171_n N_VSS_c_173_n N_VSS_c_174_n N_VSS_c_175_n
+ N_VSS_c_281_p N_VSS_c_177_n N_VSS_c_242_p N_VSS_c_178_n N_VSS_c_183_n
+ N_VSS_c_186_n N_VSS_c_190_n N_VSS_c_194_n N_VSS_c_197_n N_VSS_c_198_n
+ N_VSS_c_201_n N_VSS_c_205_n N_VSS_c_209_n N_VSS_c_212_n N_VSS_c_214_n
+ N_VSS_c_215_n N_VSS_c_216_n N_VSS_c_220_n N_VSS_c_221_n VSS N_VSS_c_226_n
+ N_VSS_c_227_n N_VSS_c_228_n Vss PM_G5_XNOR3_N3_VSS
x_PM_G5_XNOR3_N3_CI N_CI_XI22.X0_D N_CI_XI26.X0_D N_CI_XI27.X0_S N_CI_XI28.X0_S
+ N_CI_c_285_n N_CI_c_297_n N_CI_c_326_p N_CI_c_286_n N_CI_c_304_n N_CI_c_328_p
+ N_CI_c_290_n N_CI_c_310_n N_CI_c_313_p N_CI_c_322_p Vss PM_G5_XNOR3_N3_CI
x_PM_G5_XNOR3_N3_A N_A_XI21.X0_CG N_A_XI24.X0_CG N_A_XI29.X0_PGD N_A_XI28.X0_PGD
+ N_A_c_332_n N_A_c_361_p N_A_c_373_p N_A_c_375_p N_A_c_333_n N_A_c_338_n
+ N_A_c_339_n N_A_c_340_n A N_A_c_346_n N_A_c_347_n N_A_c_341_n N_A_c_364_p Vss
+ PM_G5_XNOR3_N3_A
x_PM_G5_XNOR3_N3_BI N_BI_XI25.X0_D N_BI_XI23.X0_D N_BI_XI27.X0_CG
+ N_BI_XI29.X0_CG N_BI_c_432_p N_BI_c_423_n N_BI_c_401_n N_BI_c_403_n
+ N_BI_c_437_p N_BI_c_418_n N_BI_c_433_p N_BI_c_427_n N_BI_c_408_n N_BI_c_416_n
+ N_BI_c_431_n N_BI_c_409_n N_BI_c_458_p N_BI_c_410_n Vss PM_G5_XNOR3_N3_BI
x_PM_G5_XNOR3_N3_AI N_AI_XI21.X0_D N_AI_XI24.X0_D N_AI_XI31.X0_PGD
+ N_AI_XI27.X0_PGD N_AI_c_478_n N_AI_c_469_n N_AI_c_470_n N_AI_c_472_n
+ N_AI_c_476_n N_AI_c_485_n N_AI_c_486_n Vss PM_G5_XNOR3_N3_AI
x_PM_G5_XNOR3_N3_B N_B_XI25.X0_CG N_B_XI23.X0_CG N_B_XI31.X0_CG N_B_XI28.X0_CG
+ N_B_c_515_n N_B_c_516_n N_B_c_522_n N_B_c_532_n B N_B_c_535_n N_B_c_526_n
+ N_B_c_537_n N_B_c_540_n N_B_c_542_n N_B_c_517_n N_B_c_563_n N_B_c_566_n Vss
+ PM_G5_XNOR3_N3_B
x_PM_G5_XNOR3_N3_Z N_Z_XI31.X0_D N_Z_XI27.X0_D N_Z_XI29.X0_D N_Z_XI28.X0_D
+ N_Z_c_577_n N_Z_c_584_n N_Z_c_581_n Z Vss PM_G5_XNOR3_N3_Z
cc_1 N_VDD_XI25.X0_PGD N_C_XI26.X0_CG 0.00111653f
cc_2 N_VDD_c_2_p N_C_XI26.X0_CG 0.00108697f
cc_3 N_VDD_XI26.X0_PGD N_C_c_116_n 4.20258e-19
cc_4 N_VDD_c_4_p N_C_c_116_n 0.00111653f
cc_5 N_VDD_c_5_p N_C_c_116_n 0.00135138f
cc_6 N_VDD_c_6_p N_C_c_119_n 3.43419e-19
cc_7 N_VDD_c_7_p N_C_c_120_n 4.76491e-19
cc_8 N_VDD_c_5_p N_C_c_120_n 0.00161703f
cc_9 N_VDD_c_5_p N_C_c_122_n 2.84771e-19
cc_10 N_VDD_c_10_p N_C_c_123_n 5.71495e-19
cc_11 N_VDD_c_11_p N_C_c_123_n 8.59389e-19
cc_12 N_VDD_XI26.X0_PGD N_VSS_XI22.X0_PGD 0.00200994f
cc_13 N_VDD_c_13_p N_VSS_XI22.X0_PGD 4.18763e-19
cc_14 N_VDD_XI25.X0_PGD N_VSS_XI21.X0_PGD 2.44446e-19
cc_15 N_VDD_XI24.X0_PGD N_VSS_XI21.X0_PGD 0.00200236f
cc_16 N_VDD_c_16_p N_VSS_XI21.X0_PGD 4.15609e-19
cc_17 N_VDD_XI25.X0_PGD N_VSS_XI23.X0_PGD 0.00200584f
cc_18 N_VDD_XI24.X0_PGD N_VSS_XI23.X0_PGD 2.31309e-19
cc_19 N_VDD_c_19_p N_VSS_c_170_n 0.00200994f
cc_20 N_VDD_c_20_p N_VSS_c_171_n 0.00200236f
cc_21 N_VDD_c_21_p N_VSS_c_171_n 3.00203e-19
cc_22 N_VDD_c_21_p N_VSS_c_173_n 3.89167e-19
cc_23 N_VDD_c_11_p N_VSS_c_174_n 2.35465e-19
cc_24 N_VDD_c_24_p N_VSS_c_175_n 0.00200584f
cc_25 N_VDD_c_25_p N_VSS_c_175_n 3.89167e-19
cc_26 N_VDD_c_5_p N_VSS_c_177_n 2.74986e-19
cc_27 N_VDD_c_13_p N_VSS_c_178_n 4.32468e-19
cc_28 N_VDD_c_5_p N_VSS_c_178_n 3.08724e-19
cc_29 N_VDD_c_29_p N_VSS_c_178_n 0.00111881f
cc_30 N_VDD_c_30_p N_VSS_c_178_n 3.98949e-19
cc_31 N_VDD_c_2_p N_VSS_c_178_n 3.48267e-19
cc_32 N_VDD_c_5_p N_VSS_c_183_n 2.9533e-19
cc_33 N_VDD_c_10_p N_VSS_c_183_n 7.43603e-19
cc_34 N_VDD_c_11_p N_VSS_c_183_n 8.20353e-19
cc_35 N_VDD_c_16_p N_VSS_c_186_n 6.9475e-19
cc_36 N_VDD_c_21_p N_VSS_c_186_n 0.00161703f
cc_37 N_VDD_c_37_p N_VSS_c_186_n 9.10421e-19
cc_38 N_VDD_c_38_p N_VSS_c_186_n 3.48267e-19
cc_39 N_VDD_c_10_p N_VSS_c_190_n 4.06132e-19
cc_40 N_VDD_c_25_p N_VSS_c_190_n 0.00161703f
cc_41 N_VDD_c_11_p N_VSS_c_190_n 0.00146019f
cc_42 N_VDD_c_42_p N_VSS_c_190_n 3.48267e-19
cc_43 N_VDD_XI24.X0_PGD N_VSS_c_194_n 2.99706e-19
cc_44 N_VDD_c_37_p N_VSS_c_194_n 0.00524008f
cc_45 N_VDD_c_38_p N_VSS_c_194_n 9.58524e-19
cc_46 N_VDD_c_21_p N_VSS_c_197_n 0.00400652f
cc_47 N_VDD_c_13_p N_VSS_c_198_n 4.41003e-19
cc_48 N_VDD_c_30_p N_VSS_c_198_n 3.89161e-19
cc_49 N_VDD_c_2_p N_VSS_c_198_n 7.99831e-19
cc_50 N_VDD_c_16_p N_VSS_c_201_n 3.48267e-19
cc_51 N_VDD_c_21_p N_VSS_c_201_n 2.26455e-19
cc_52 N_VDD_c_37_p N_VSS_c_201_n 3.99794e-19
cc_53 N_VDD_c_38_p N_VSS_c_201_n 6.489e-19
cc_54 N_VDD_c_10_p N_VSS_c_205_n 3.82294e-19
cc_55 N_VDD_c_25_p N_VSS_c_205_n 2.26455e-19
cc_56 N_VDD_c_11_p N_VSS_c_205_n 9.55109e-19
cc_57 N_VDD_c_42_p N_VSS_c_205_n 6.46219e-19
cc_58 N_VDD_c_7_p N_VSS_c_209_n 0.00419405f
cc_59 N_VDD_c_13_p N_VSS_c_209_n 0.00325114f
cc_60 N_VDD_c_60_p N_VSS_c_209_n 0.0010705f
cc_61 N_VDD_c_13_p N_VSS_c_212_n 0.0102114f
cc_62 N_VDD_c_30_p N_VSS_c_212_n 0.00124944f
cc_63 N_VDD_c_5_p N_VSS_c_214_n 0.0097003f
cc_64 N_VDD_c_64_p N_VSS_c_215_n 0.00107633f
cc_65 N_VDD_c_65_p N_VSS_c_216_n 0.00833289f
cc_66 N_VDD_c_66_p N_VSS_c_216_n 6.51257e-19
cc_67 N_VDD_c_21_p N_VSS_c_216_n 0.00369311f
cc_68 N_VDD_c_68_p N_VSS_c_216_n 0.00146091f
cc_69 N_VDD_c_69_p N_VSS_c_220_n 0.00107845f
cc_70 N_VDD_c_5_p N_VSS_c_221_n 0.00143483f
cc_71 N_VDD_c_25_p N_VSS_c_221_n 0.00610315f
cc_72 N_VDD_c_72_p N_VSS_c_221_n 9.53204e-19
cc_73 N_VDD_c_10_p VSS 2.72347e-19
cc_74 N_VDD_c_11_p VSS 9.64592e-19
cc_75 N_VDD_c_13_p N_VSS_c_226_n 0.00109802f
cc_76 N_VDD_c_5_p N_VSS_c_227_n 0.00111918f
cc_77 N_VDD_c_21_p N_VSS_c_228_n 7.74609e-19
cc_78 N_VDD_c_78_p N_CI_c_285_n 3.43419e-19
cc_79 N_VDD_c_78_p N_CI_c_286_n 3.48267e-19
cc_80 N_VDD_c_5_p N_CI_c_286_n 3.21336e-19
cc_81 N_VDD_c_29_p N_CI_c_286_n 5.61123e-19
cc_82 N_VDD_c_30_p N_CI_c_286_n 0.00278407f
cc_83 N_VDD_c_16_p N_CI_c_290_n 7.63838e-19
cc_84 N_VDD_c_66_p N_CI_c_290_n 4.68699e-19
cc_85 N_VDD_XI24.X0_PGD N_A_c_332_n 3.96972e-19
cc_86 N_VDD_XI24.X0_PGD N_A_c_333_n 5.06189e-19
cc_87 N_VDD_c_6_p N_A_c_333_n 2.21087e-19
cc_88 N_VDD_c_21_p N_A_c_333_n 2.0692e-19
cc_89 N_VDD_c_11_p N_A_c_333_n 3.17218e-19
cc_90 N_VDD_c_38_p N_A_c_333_n 2.03128e-19
cc_91 N_VDD_c_6_p N_A_c_338_n 9.18655e-19
cc_92 N_VDD_c_11_p N_A_c_339_n 0.0068268f
cc_93 N_VDD_c_30_p N_A_c_340_n 0.00109781f
cc_94 N_VDD_c_30_p N_A_c_341_n 5.7233e-19
cc_95 N_VDD_c_6_p N_BI_c_401_n 3.43419e-19
cc_96 N_VDD_c_11_p N_BI_c_401_n 3.48267e-19
cc_97 N_VDD_c_6_p N_BI_c_403_n 3.48267e-19
cc_98 N_VDD_c_30_p N_BI_c_403_n 7.69656e-19
cc_99 N_VDD_c_25_p N_BI_c_403_n 3.21336e-19
cc_100 N_VDD_c_11_p N_BI_c_403_n 4.99861e-19
cc_101 N_VDD_XI24.X0_PGD N_AI_XI31.X0_PGD 3.10667e-19
cc_102 N_VDD_c_102_p N_AI_c_469_n 3.10667e-19
cc_103 N_VDD_c_103_p N_AI_c_470_n 3.43419e-19
cc_104 N_VDD_c_66_p N_AI_c_470_n 3.73302e-19
cc_105 N_VDD_c_103_p N_AI_c_472_n 3.48267e-19
cc_106 N_VDD_c_16_p N_AI_c_472_n 3.47482e-19
cc_107 N_VDD_c_66_p N_AI_c_472_n 5.23123e-19
cc_108 N_VDD_c_21_p N_AI_c_472_n 3.21336e-19
cc_109 N_VDD_c_37_p N_AI_c_476_n 0.00118673f
cc_110 N_VDD_XI26.X0_PGD N_B_XI25.X0_CG 0.00111782f
cc_111 N_VDD_XI25.X0_PGD N_B_c_515_n 4.01605e-19
cc_112 N_VDD_c_112_p N_B_c_516_n 0.00111782f
cc_113 N_VDD_c_11_p N_B_c_517_n 4.72333e-19
cc_114 N_C_c_116_n N_VSS_XI22.X0_PGD 4.20258e-19
cc_115 N_C_c_126_p N_VSS_c_230_n 2.76939e-19
cc_116 N_C_c_127_p N_VSS_c_183_n 7.31268e-19
cc_117 N_C_c_123_n N_VSS_c_183_n 0.00200258f
cc_118 N_C_c_129_p N_VSS_c_198_n 0.0041528f
cc_119 N_C_c_120_n N_VSS_c_209_n 4.01014e-19
cc_120 N_C_c_123_n N_VSS_c_209_n 2.67373e-19
cc_121 N_C_c_120_n N_VSS_c_214_n 0.00171716f
cc_122 N_C_c_123_n N_VSS_c_214_n 0.00318423f
cc_123 N_C_c_123_n N_VSS_c_221_n 0.00192963f
cc_124 N_C_c_123_n VSS 0.00167449f
cc_125 N_C_c_116_n N_CI_c_285_n 7.69306e-19
cc_126 N_C_c_123_n N_CI_c_286_n 7.42955e-19
cc_127 N_C_c_123_n N_CI_c_290_n 0.00148047f
cc_128 N_C_c_123_n N_A_c_333_n 3.38948e-19
cc_129 N_C_c_119_n N_A_c_338_n 8.20481e-19
cc_130 N_C_c_127_p N_A_c_338_n 0.00202163f
cc_131 N_C_c_123_n N_A_c_339_n 5.50651e-19
cc_132 N_C_c_143_p N_A_c_346_n 7.67297e-19
cc_133 N_C_c_119_n N_A_c_347_n 5.83331e-19
cc_134 N_C_c_127_p N_A_c_347_n 0.00118769f
cc_135 N_C_c_123_n N_A_c_347_n 4.69432e-19
cc_136 N_C_c_143_p N_A_c_347_n 0.00239654f
cc_137 N_C_c_148_p N_A_c_347_n 3.74525e-19
cc_138 N_C_c_123_n N_BI_c_403_n 2.74336e-19
cc_139 N_C_c_123_n N_BI_c_408_n 3.41448e-19
cc_140 N_C_c_143_p N_BI_c_409_n 4.45126e-19
cc_141 N_C_c_143_p N_BI_c_410_n 0.00127751f
cc_142 N_C_c_127_p N_B_c_517_n 0.00140507f
cc_143 N_C_c_123_n N_B_c_517_n 0.00214978f
cc_144 N_C_c_143_p N_B_c_517_n 9.13922e-19
cc_145 N_C_c_119_n N_Z_c_577_n 3.43419e-19
cc_146 N_C_c_157_p N_Z_c_577_n 3.43419e-19
cc_147 N_C_c_127_p N_Z_c_577_n 3.48267e-19
cc_148 N_C_c_159_p N_Z_c_577_n 3.48267e-19
cc_149 N_C_c_157_p N_Z_c_581_n 3.48267e-19
cc_150 N_C_c_127_p N_Z_c_581_n 6.09821e-19
cc_151 N_C_c_159_p N_Z_c_581_n 5.71987e-19
cc_152 N_VSS_c_177_n N_CI_c_285_n 3.43419e-19
cc_153 N_VSS_c_183_n N_CI_c_285_n 3.48267e-19
cc_154 N_VSS_c_242_p N_CI_c_297_n 3.43419e-19
cc_155 N_VSS_c_194_n N_CI_c_297_n 3.48267e-19
cc_156 N_VSS_c_177_n N_CI_c_286_n 3.48267e-19
cc_157 N_VSS_c_178_n N_CI_c_286_n 5.78167e-19
cc_158 N_VSS_c_183_n N_CI_c_286_n 0.00107566f
cc_159 N_VSS_c_209_n N_CI_c_286_n 6.53442e-19
cc_160 N_VSS_c_212_n N_CI_c_286_n 0.00285518f
cc_161 N_VSS_c_242_p N_CI_c_304_n 3.48267e-19
cc_162 N_VSS_c_194_n N_CI_c_304_n 0.00120696f
cc_163 N_VSS_c_186_n N_CI_c_290_n 0.00138401f
cc_164 N_VSS_c_194_n N_CI_c_290_n 2.05251e-19
cc_165 N_VSS_c_197_n N_CI_c_290_n 0.00334374f
cc_166 N_VSS_c_216_n N_CI_c_290_n 2.16087e-19
cc_167 N_VSS_c_216_n N_CI_c_310_n 0.00293637f
cc_168 N_VSS_XI21.X0_PGD N_A_c_332_n 3.96972e-19
cc_169 N_VSS_c_242_p N_A_c_333_n 4.13509e-19
cc_170 N_VSS_c_194_n N_A_c_333_n 7.30817e-19
cc_171 N_VSS_c_197_n N_A_c_333_n 2.62883e-19
cc_172 N_VSS_c_201_n N_A_c_340_n 2.09367e-19
cc_173 N_VSS_c_186_n N_A_c_341_n 2.04211e-19
cc_174 N_VSS_c_201_n N_A_c_341_n 4.89964e-19
cc_175 N_VSS_c_177_n N_BI_c_401_n 3.43419e-19
cc_176 N_VSS_c_183_n N_BI_c_401_n 3.48267e-19
cc_177 N_VSS_c_177_n N_BI_c_403_n 3.48267e-19
cc_178 N_VSS_c_183_n N_BI_c_403_n 0.00101872f
cc_179 N_VSS_c_221_n N_BI_c_403_n 2.19864e-19
cc_180 N_VSS_c_197_n N_BI_c_416_n 2.2551e-19
cc_181 N_VSS_XI23.X0_PGD N_AI_XI31.X0_PGD 2.79882e-19
cc_182 N_VSS_c_174_n N_AI_c_478_n 2.79882e-19
cc_183 N_VSS_c_242_p N_AI_c_470_n 3.43419e-19
cc_184 N_VSS_c_194_n N_AI_c_470_n 3.48267e-19
cc_185 N_VSS_c_242_p N_AI_c_472_n 3.48267e-19
cc_186 N_VSS_c_194_n N_AI_c_472_n 0.00173694f
cc_187 N_VSS_c_194_n N_AI_c_476_n 0.00177896f
cc_188 N_VSS_c_197_n N_AI_c_476_n 0.00605709f
cc_189 N_VSS_c_194_n N_AI_c_485_n 2.82216e-19
cc_190 N_VSS_c_186_n N_AI_c_486_n 0.00195338f
cc_191 N_VSS_c_197_n N_AI_c_486_n 0.00167789f
cc_192 N_VSS_XI23.X0_PGD N_B_c_515_n 4.01605e-19
cc_193 N_VSS_c_281_p N_B_c_522_n 6.24637e-19
cc_194 N_VSS_c_190_n B 2.2661e-19
cc_195 N_VSS_c_205_n B 2.39151e-19
cc_196 VSS N_B_c_517_n 2.35905e-19
cc_197 N_CI_c_290_n N_A_c_333_n 3.7003e-19
cc_198 N_CI_c_286_n N_BI_c_403_n 0.00144806f
cc_199 N_CI_c_313_p N_BI_c_418_n 5.10764e-19
cc_200 N_CI_c_304_n N_BI_c_408_n 6.46554e-19
cc_201 N_CI_c_290_n N_BI_c_408_n 8.14649e-19
cc_202 N_CI_c_313_p N_BI_c_409_n 0.0012701f
cc_203 N_CI_c_286_n N_AI_c_472_n 8.00553e-19
cc_204 N_CI_c_304_n N_AI_c_472_n 9.98055e-19
cc_205 N_CI_c_304_n N_AI_c_476_n 0.00117248f
cc_206 N_CI_c_290_n N_AI_c_476_n 0.00763297f
cc_207 N_CI_c_313_p N_AI_c_476_n 0.00313643f
cc_208 N_CI_c_322_p N_AI_c_476_n 0.00100316f
cc_209 N_CI_c_290_n N_AI_c_486_n 9.91646e-19
cc_210 N_CI_c_313_p N_B_c_526_n 7.08144e-19
cc_211 N_CI_c_297_n N_Z_c_584_n 3.43419e-19
cc_212 N_CI_c_326_p N_Z_c_584_n 3.43419e-19
cc_213 N_CI_c_304_n N_Z_c_584_n 3.48267e-19
cc_214 N_CI_c_328_p N_Z_c_584_n 3.48267e-19
cc_215 N_CI_c_326_p N_Z_c_581_n 3.48267e-19
cc_216 N_CI_c_304_n N_Z_c_581_n 6.09821e-19
cc_217 N_CI_c_328_p N_Z_c_581_n 5.71987e-19
cc_218 N_A_XI29.X0_PGD N_BI_XI29.X0_CG 9.65637e-19
cc_219 N_A_c_361_p N_BI_c_423_n 5.35095e-19
cc_220 N_A_c_333_n N_BI_c_403_n 3.00325e-19
cc_221 N_A_c_338_n N_BI_c_403_n 0.00110499f
cc_222 N_A_c_364_p N_BI_c_418_n 2.15082e-19
cc_223 N_A_XI29.X0_PGD N_BI_c_427_n 0.00133285f
cc_224 N_A_c_346_n N_BI_c_427_n 2.15082e-19
cc_225 N_A_c_338_n N_BI_c_408_n 0.00187419f
cc_226 N_A_c_333_n N_BI_c_416_n 0.00339867f
cc_227 N_A_c_338_n N_BI_c_431_n 3.69994e-19
cc_228 N_A_XI29.X0_PGD N_AI_XI31.X0_PGD 0.0173493f
cc_229 N_A_c_338_n N_AI_XI31.X0_PGD 0.001002f
cc_230 N_A_c_347_n N_AI_XI31.X0_PGD 7.67512e-19
cc_231 N_A_c_373_p N_AI_c_478_n 0.00199603f
cc_232 N_A_c_347_n N_AI_c_478_n 0.00128901f
cc_233 N_A_c_375_p N_AI_c_469_n 0.00201004f
cc_234 N_A_c_332_n N_AI_c_470_n 6.90199e-19
cc_235 N_A_c_333_n N_AI_c_472_n 5.84011e-19
cc_236 N_A_c_333_n N_AI_c_476_n 0.00127614f
cc_237 N_A_c_332_n N_B_c_515_n 0.00360349f
cc_238 N_A_c_333_n N_B_c_515_n 5.25071e-19
cc_239 N_A_c_340_n N_B_c_516_n 5.25071e-19
cc_240 N_A_c_341_n N_B_c_516_n 7.41063e-19
cc_241 N_A_c_333_n N_B_c_522_n 3.90215e-19
cc_242 N_A_XI29.X0_PGD N_B_c_532_n 9.65637e-19
cc_243 N_A_c_333_n B 6.34584e-19
cc_244 N_A_c_338_n B 4.3123e-19
cc_245 N_A_c_338_n N_B_c_535_n 4.01937e-19
cc_246 N_A_c_347_n N_B_c_535_n 3.79361e-19
cc_247 N_A_c_332_n N_B_c_537_n 7.73422e-19
cc_248 N_A_c_333_n N_B_c_537_n 5.77217e-19
cc_249 N_A_c_338_n N_B_c_537_n 6.37149e-19
cc_250 N_A_c_338_n N_B_c_540_n 3.37713e-19
cc_251 N_A_c_347_n N_B_c_540_n 2.21087e-19
cc_252 N_A_XI29.X0_PGD N_B_c_542_n 0.00133285f
cc_253 N_A_c_338_n N_B_c_517_n 0.00197838f
cc_254 N_A_c_347_n N_B_c_517_n 0.00180845f
cc_255 N_A_c_347_n N_Z_c_577_n 7.79328e-19
cc_256 N_A_XI29.X0_PGD N_Z_c_581_n 7.77706e-19
cc_257 N_A_c_338_n N_Z_c_581_n 0.00169143f
cc_258 N_A_c_347_n N_Z_c_581_n 0.0010247f
cc_259 N_BI_c_432_p N_AI_XI31.X0_PGD 9.65637e-19
cc_260 N_BI_c_433_p N_AI_XI31.X0_PGD 0.00133285f
cc_261 N_BI_c_416_n N_AI_c_472_n 6.07277e-19
cc_262 N_BI_c_433_p N_AI_c_476_n 2.15082e-19
cc_263 N_BI_c_408_n N_AI_c_476_n 0.00233431f
cc_264 N_BI_c_437_p N_AI_c_485_n 2.15082e-19
cc_265 N_BI_c_433_p N_AI_c_485_n 5.05931e-19
cc_266 N_BI_c_401_n N_B_c_515_n 6.90199e-19
cc_267 N_BI_c_403_n B 5.19468e-19
cc_268 N_BI_c_408_n B 2.66639e-19
cc_269 N_BI_c_437_p N_B_c_535_n 3.94971e-19
cc_270 N_BI_c_433_p N_B_c_535_n 4.03665e-19
cc_271 N_BI_c_408_n N_B_c_535_n 2.81186e-19
cc_272 N_BI_c_418_n N_B_c_526_n 0.00181951f
cc_273 N_BI_c_427_n N_B_c_526_n 4.56568e-19
cc_274 N_BI_c_437_p N_B_c_540_n 4.44913e-19
cc_275 N_BI_c_433_p N_B_c_540_n 0.00360065f
cc_276 N_BI_c_427_n N_B_c_540_n 0.00102603f
cc_277 N_BI_c_433_p N_B_c_542_n 7.16621e-19
cc_278 N_BI_c_427_n N_B_c_542_n 0.00243716f
cc_279 N_BI_c_403_n N_B_c_517_n 0.00150424f
cc_280 N_BI_c_418_n N_B_c_517_n 0.00163797f
cc_281 N_BI_c_408_n N_B_c_517_n 0.0161531f
cc_282 N_BI_c_409_n N_B_c_517_n 8.58649e-19
cc_283 N_BI_c_410_n N_B_c_517_n 6.57534e-19
cc_284 N_BI_c_408_n N_B_c_563_n 0.0022474f
cc_285 N_BI_c_458_p N_B_c_563_n 0.00206348f
cc_286 N_BI_c_410_n N_B_c_563_n 2.41136e-19
cc_287 N_BI_c_437_p N_B_c_566_n 3.09421e-19
cc_288 N_BI_c_431_n N_B_c_566_n 0.0022474f
cc_289 N_BI_c_409_n N_B_c_566_n 8.20948e-19
cc_290 N_BI_c_437_p N_Z_c_581_n 0.00157325f
cc_291 N_BI_c_418_n N_Z_c_581_n 0.00155051f
cc_292 N_BI_c_433_p N_Z_c_581_n 8.66889e-19
cc_293 N_BI_c_427_n N_Z_c_581_n 8.66889e-19
cc_294 N_BI_c_408_n N_Z_c_581_n 3.95297e-19
cc_295 N_AI_XI31.X0_PGD N_B_XI31.X0_CG 9.47088e-19
cc_296 N_AI_XI31.X0_PGD N_B_c_540_n 0.00340539f
cc_297 N_AI_XI31.X0_PGD N_Z_c_581_n 4.24987e-19
cc_298 N_B_c_535_n N_Z_c_581_n 0.00158441f
cc_299 N_B_c_526_n N_Z_c_581_n 0.00138952f
cc_300 N_B_c_542_n N_Z_c_581_n 8.66889e-19
cc_301 N_B_c_517_n N_Z_c_581_n 7.81804e-19
cc_302 N_B_c_563_n N_Z_c_581_n 0.00232585f
cc_303 N_B_c_566_n N_Z_c_581_n 0.00104129f
*
.ends
*
*
.subckt XNOR3_HPNW12 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XNOR3_N3
.ends
*
* File: G4_XOR2_N3.pex.netlist
* Created: Sun Apr 10 19:09:34 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XOR2_N3_VSS 2 5 9 12 14 16 32 33 42 43 54 59 63 66 71 76 81 86 95
+ 100 113 115 116 117 122 123 128 138 140 145 146 147 150 Vss
c92 148 Vss 6.20041e-19
c93 147 Vss 3.75522e-19
c94 146 Vss 4.28045e-19
c95 145 Vss 0.00444873f
c96 140 Vss 0.00219072f
c97 138 Vss 0.00853623f
c98 128 Vss 0.00370986f
c99 123 Vss 8.46757e-19
c100 122 Vss 0.00174135f
c101 117 Vss 8.2479e-19
c102 116 Vss 0.00447709f
c103 115 Vss 0.00650684f
c104 113 Vss 0.00239513f
c105 100 Vss 0.00529998f
c106 95 Vss 0.00418654f
c107 86 Vss 2.86598e-19
c108 81 Vss 0.00160268f
c109 76 Vss 0.0010261f
c110 71 Vss 0.00123398f
c111 66 Vss 0.00174721f
c112 63 Vss 0.0101876f
c113 59 Vss 0.00691967f
c114 54 Vss 0.0100924f
c115 43 Vss 0.0342915f
c116 42 Vss 0.100071f
c117 33 Vss 0.0350852f
c118 32 Vss 0.0990727f
c119 14 Vss 0.00143493f
c120 9 Vss 0.384391f
c121 5 Vss 0.378692f
r122 145 150 0.326018
r123 144 145 5.50157
r124 140 144 0.655813
r125 139 148 0.494161
r126 138 150 0.326018
r127 138 139 13.0037
r128 134 148 0.128424
r129 129 147 0.494161
r130 128 148 0.494161
r131 128 129 7.46046
r132 124 147 0.128424
r133 122 147 0.494161
r134 122 123 4.37625
r135 118 146 0.0828784
r136 116 130 0.652036
r137 116 117 10.1279
r138 115 123 0.652036
r139 114 146 0.551426
r140 114 115 17.1716
r141 113 146 0.551426
r142 112 117 0.652036
r143 112 113 5.79332
r144 86 140 1.82344
r145 81 134 6.16843
r146 76 100 1.16709
r147 76 130 2.16729
r148 71 95 1.16709
r149 71 124 2.16729
r150 66 118 1.82344
r151 63 86 1.16709
r152 59 81 1.16709
r153 54 66 1.16709
r154 45 100 0.119107
r155 43 45 1.45875
r156 42 46 0.652036
r157 42 45 1.45875
r158 39 43 0.652036
r159 35 95 0.0476429
r160 33 35 1.45875
r161 32 36 0.652036
r162 32 35 1.45875
r163 29 33 0.652036
r164 16 63 0.123773
r165 14 59 0.123773
r166 12 59 0.123773
r167 9 46 5.1348
r168 9 39 5.1348
r169 5 36 5.1348
r170 5 29 5.1348
r171 2 54 0.123773
.ends

.subckt PM_G4_XOR2_N3_VDD 3 6 8 11 14 16 32 42 43 54 59 66 68 69 70 73 75 76 79
+ 81 85 89 91 93 98 99 100 103 109 114 123 Vss
c98 123 Vss 0.00813195f
c99 114 Vss 0.00444328f
c100 109 Vss 0.00562387f
c101 101 Vss 8.87755e-19
c102 100 Vss 2.39889e-19
c103 99 Vss 4.52364e-19
c104 98 Vss 0.0063791f
c105 93 Vss 0.00162315f
c106 91 Vss 0.0131786f
c107 89 Vss 0.00230903f
c108 85 Vss 7.1324e-19
c109 81 Vss 0.00459876f
c110 79 Vss 0.00140429f
c111 76 Vss 8.64616e-19
c112 75 Vss 0.00587269f
c113 73 Vss 0.00191373f
c114 70 Vss 8.68689e-19
c115 69 Vss 0.00224797f
c116 68 Vss 0.00279777f
c117 66 Vss 0.0108403f
c118 59 Vss 0.00695462f
c119 54 Vss 0.00822951f
c120 43 Vss 0.0351405f
c121 42 Vss 0.100972f
c122 33 Vss 0.0359366f
c123 32 Vss 0.100971f
c124 14 Vss 0.00143493f
c125 11 Vss 0.377105f
c126 3 Vss 0.384936f
r127 98 103 0.349767
r128 97 98 5.75164
r129 95 123 1.16709
r130 93 103 0.306046
r131 93 95 1.82344
r132 92 101 0.494161
r133 91 97 0.652036
r134 91 92 13.0037
r135 87 101 0.128424
r136 87 89 6.46018
r137 85 114 1.16709
r138 83 85 2.16729
r139 82 100 0.494161
r140 81 101 0.494161
r141 81 82 7.46046
r142 79 109 1.16709
r143 77 100 0.128424
r144 77 79 2.16729
r145 75 83 0.652036
r146 75 76 10.1279
r147 71 99 0.0828784
r148 71 73 1.82344
r149 69 100 0.494161
r150 69 70 4.37625
r151 68 76 0.652036
r152 67 99 0.551426
r153 67 68 5.50157
r154 66 99 0.551426
r155 65 70 0.652036
r156 65 66 17.4633
r157 63 123 0.05
r158 59 89 1.16709
r159 54 73 1.02121
r160 45 114 0.0476429
r161 43 45 1.45875
r162 42 46 0.652036
r163 42 45 1.45875
r164 39 43 0.652036
r165 35 109 0.119107
r166 33 35 1.45875
r167 32 36 0.652036
r168 32 35 1.45875
r169 29 33 0.652036
r170 16 63 0.123773
r171 14 59 0.123773
r172 11 46 5.1348
r173 11 39 5.1348
r174 8 59 0.123773
r175 6 54 0.123773
r176 3 36 5.1348
r177 3 29 5.1348
.ends

.subckt PM_G4_XOR2_N3_A 2 4 7 10 21 24 28 48 51 54 57 62 67 72 77 85 Vss
c54 85 Vss 8.24403e-19
c55 77 Vss 0.00191043f
c56 72 Vss 0.00680655f
c57 67 Vss 0.00366581f
c58 62 Vss 0.00280314f
c59 57 Vss 0.00457389f
c60 51 Vss 0.00108099f
c61 48 Vss 0.128068f
c62 43 Vss 0.0296639f
c63 28 Vss 0.152693f
c64 24 Vss 8.47557e-20
c65 21 Vss 0.173351f
c66 18 Vss 0.180502f
c67 16 Vss 0.0247918f
c68 10 Vss 0.176342f
c69 7 Vss 0.432086f
c70 4 Vss 0.193054f
r71 81 85 0.653045
r72 62 77 1.16709
r73 62 85 4.9014
r74 57 72 1.16709
r75 57 81 10.8364
r76 51 67 1.16709
r77 51 54 0.0833571
r78 47 72 0.0238214
r79 47 48 2.334
r80 44 47 2.20433
r81 39 77 0.50025
r82 33 48 0.00605528
r83 31 44 0.00605528
r84 29 43 0.494161
r85 28 30 0.652036
r86 28 29 4.84305
r87 25 43 0.128424
r88 24 67 0.0476429
r89 22 24 0.326018
r90 22 24 0.1167
r91 21 43 0.494161
r92 21 24 6.7686
r93 18 67 0.357321
r94 16 24 0.326018
r95 16 18 0.40845
r96 10 39 4.668
r97 7 33 5.1348
r98 7 31 5.1348
r99 7 30 5.1348
r100 4 25 5.1348
r101 2 18 4.72635
.ends

.subckt PM_G4_XOR2_N3_NET1 2 4 7 10 31 35 41 44 49 58 76 Vss
c34 76 Vss 3.97901e-19
c35 58 Vss 0.0058132f
c36 49 Vss 0.00651255f
c37 44 Vss 0.00236298f
c38 41 Vss 0.00514975f
c39 35 Vss 0.103147f
c40 31 Vss 0.12549f
c41 10 Vss 0.269166f
c42 7 Vss 0.499657f
c43 4 Vss 0.00143493f
r44 72 76 0.655813
r45 49 58 1.16709
r46 49 76 12.1076
r47 44 72 3.62604
r48 41 44 1.16709
r49 33 35 1.70187
r50 30 58 0.142929
r51 30 31 2.20433
r52 27 30 2.334
r53 25 35 0.17282
r54 24 31 0.00605528
r55 21 33 0.17282
r56 18 27 0.00605528
r57 10 21 7.64385
r58 7 25 7.29375
r59 7 24 5.1348
r60 7 18 5.1348
r61 4 41 0.123773
r62 2 41 0.123773
.ends

.subckt PM_G4_XOR2_N3_NET2 2 4 6 9 21 22 33 39 42 47 56 74 Vss
c42 74 Vss 3.21991e-19
c43 56 Vss 0.00502059f
c44 47 Vss 0.00781175f
c45 42 Vss 0.00242715f
c46 39 Vss 0.00509494f
c47 33 Vss 0.12909f
c48 22 Vss 0.0345713f
c49 21 Vss 0.177367f
c50 9 Vss 0.573605f
c51 6 Vss 0.188648f
c52 4 Vss 0.00143493f
r53 70 74 0.660011
r54 47 56 1.16709
r55 47 74 11.3611
r56 42 70 3.29261
r57 39 42 1.16709
r58 32 56 0.0238214
r59 32 33 2.26917
r60 29 32 2.26917
r61 26 33 0.00605528
r62 24 29 0.00605528
r63 21 23 0.652036
r64 21 22 4.84305
r65 18 22 0.652036
r66 9 26 5.1348
r67 9 24 5.1348
r68 9 23 10.0362
r69 6 18 5.1348
r70 4 39 0.123773
r71 2 39 0.123773
.ends

.subckt PM_G4_XOR2_N3_B 2 4 7 10 19 20 28 31 35 45 51 54 Vss
c31 54 Vss 0.0283542f
c32 51 Vss 0.00177471f
c33 45 Vss 0.13328f
c34 35 Vss 0.154928f
c35 31 Vss 2.04877e-19
c36 28 Vss 0.117534f
c37 20 Vss 0.0348422f
c38 19 Vss 0.173065f
c39 10 Vss 0.264298f
c40 7 Vss 0.440555f
c41 4 Vss 0.189408f
c42 2 Vss 0.201403f
r43 51 54 1.16709
r44 43 45 4.53833
r45 38 45 0.00605528
r46 35 47 1.87725
r47 33 47 0.527901
r48 32 43 0.00605528
r49 31 54 0.181909
r50 29 54 0.494161
r51 29 31 0.1167
r52 28 47 0.333556
r53 28 31 4.72635
r54 23 54 0.128424
r55 23 54 0.40845
r56 22 54 0.181909
r57 20 22 6.7686
r58 19 54 0.494161
r59 19 22 0.1167
r60 16 20 0.652036
r61 10 35 7.5855
r62 7 38 5.1348
r63 7 33 5.42655
r64 7 32 5.1348
r65 4 54 5.0181
r66 2 16 5.42655
.ends

.subckt PM_G4_XOR2_N3_Z 2 4 6 8 23 27 30 33 Vss
c29 30 Vss 0.00322833f
c30 27 Vss 0.00675283f
c31 23 Vss 0.00497092f
c32 8 Vss 0.00143493f
c33 6 Vss 0.00143493f
r34 33 35 4.95975
r35 30 33 6.71025
r36 27 35 1.16709
r37 23 30 1.16709
r38 8 27 0.123773
r39 6 23 0.123773
r40 4 27 0.123773
r41 2 23 0.123773
.ends

.subckt G4_XOR2_N3  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI20.X0 N_NET1_XI20.X0_D N_VDD_XI20.X0_PGD N_B_XI20.X0_CG N_VDD_XI20.X0_PGD
+ N_VSS_XI20.X0_S TIGFET_HPNW12
XI18.X0 N_NET2_XI18.X0_D N_VSS_XI18.X0_PGD N_A_XI18.X0_CG N_VSS_XI18.X0_PGD
+ N_VDD_XI18.X0_S TIGFET_HPNW12
XI22.X0 N_NET1_XI22.X0_D N_VSS_XI22.X0_PGD N_B_XI22.X0_CG N_VSS_XI22.X0_PGD
+ N_VDD_XI22.X0_S TIGFET_HPNW12
XI16.X0 N_NET2_XI16.X0_D N_VDD_XI16.X0_PGD N_A_XI16.X0_CG N_VDD_XI16.X0_PGD
+ N_VSS_XI16.X0_S TIGFET_HPNW12
XI21.X0 N_Z_XI21.X0_D N_B_XI21.X0_PGD N_NET2_XI21.X0_CG N_B_XI21.X0_PGD
+ N_VDD_XI21.X0_S TIGFET_HPNW12
XI19.X0 N_Z_XI19.X0_D N_A_XI19.X0_PGD N_B_XI19.X0_CG N_A_XI19.X0_PGD
+ N_VSS_XI19.X0_S TIGFET_HPNW12
XI23.X0 N_Z_XI23.X0_D N_NET1_XI23.X0_PGD N_A_XI23.X0_CG N_NET1_XI23.X0_PGD
+ N_VDD_XI23.X0_S TIGFET_HPNW12
XI17.X0 N_Z_XI17.X0_D N_NET2_XI17.X0_PGD N_NET1_XI17.X0_CG N_NET2_XI17.X0_PGD
+ N_VSS_XI17.X0_S TIGFET_HPNW12
*
x_PM_G4_XOR2_N3_VSS N_VSS_XI20.X0_S N_VSS_XI18.X0_PGD N_VSS_XI22.X0_PGD
+ N_VSS_XI16.X0_S N_VSS_XI19.X0_S N_VSS_XI17.X0_S N_VSS_c_5_p N_VSS_c_22_p
+ N_VSS_c_38_p N_VSS_c_4_p N_VSS_c_7_p N_VSS_c_6_p N_VSS_c_85_p N_VSS_c_8_p
+ N_VSS_c_13_p N_VSS_c_29_p N_VSS_c_36_p N_VSS_c_87_p N_VSS_c_14_p N_VSS_c_30_p
+ N_VSS_c_9_p N_VSS_c_10_p N_VSS_c_18_p N_VSS_c_19_p N_VSS_c_25_p N_VSS_c_28_p
+ N_VSS_c_26_p N_VSS_c_55_p N_VSS_c_41_p N_VSS_c_57_p N_VSS_c_11_p N_VSS_c_27_p
+ VSS Vss PM_G4_XOR2_N3_VSS
x_PM_G4_XOR2_N3_VDD N_VDD_XI20.X0_PGD N_VDD_XI18.X0_S N_VDD_XI22.X0_S
+ N_VDD_XI16.X0_PGD N_VDD_XI21.X0_S N_VDD_XI23.X0_S N_VDD_c_96_n N_VDD_c_144_p
+ N_VDD_c_97_n N_VDD_c_167_p N_VDD_c_98_n N_VDD_c_99_n N_VDD_c_104_n
+ N_VDD_c_108_n N_VDD_c_111_n N_VDD_c_112_n N_VDD_c_113_n N_VDD_c_120_n
+ N_VDD_c_121_n N_VDD_c_123_n N_VDD_c_127_n N_VDD_c_130_n N_VDD_c_148_p
+ N_VDD_c_133_n N_VDD_c_155_p N_VDD_c_134_n N_VDD_c_135_n VDD N_VDD_c_136_n
+ N_VDD_c_138_n N_VDD_c_185_p Vss PM_G4_XOR2_N3_VDD
x_PM_G4_XOR2_N3_A N_A_XI18.X0_CG N_A_XI16.X0_CG N_A_XI19.X0_PGD N_A_XI23.X0_CG
+ N_A_c_191_n N_A_c_193_n N_A_c_194_n N_A_c_208_n N_A_c_195_n A N_A_c_196_n
+ N_A_c_201_n N_A_c_202_n N_A_c_215_n N_A_c_219_p N_A_c_203_n Vss
+ PM_G4_XOR2_N3_A
x_PM_G4_XOR2_N3_NET1 N_NET1_XI20.X0_D N_NET1_XI22.X0_D N_NET1_XI23.X0_PGD
+ N_NET1_XI17.X0_CG N_NET1_c_250_n N_NET1_c_270_p N_NET1_c_245_n N_NET1_c_246_n
+ N_NET1_c_247_n N_NET1_c_259_n N_NET1_c_248_n Vss PM_G4_XOR2_N3_NET1
x_PM_G4_XOR2_N3_NET2 N_NET2_XI18.X0_D N_NET2_XI16.X0_D N_NET2_XI21.X0_CG
+ N_NET2_XI17.X0_PGD N_NET2_c_300_n N_NET2_c_315_p N_NET2_c_301_n N_NET2_c_279_n
+ N_NET2_c_281_n N_NET2_c_284_n N_NET2_c_306_n N_NET2_c_288_n Vss
+ PM_G4_XOR2_N3_NET2
x_PM_G4_XOR2_N3_B N_B_XI20.X0_CG N_B_XI22.X0_CG N_B_XI21.X0_PGD N_B_XI19.X0_CG
+ N_B_c_323_n N_B_c_338_n N_B_c_325_n N_B_c_326_n N_B_c_340_n N_B_c_327_n B
+ N_B_c_335_n Vss PM_G4_XOR2_N3_B
x_PM_G4_XOR2_N3_Z N_Z_XI21.X0_D N_Z_XI19.X0_D N_Z_XI23.X0_D N_Z_XI17.X0_D
+ N_Z_c_361_n N_Z_c_352_n N_Z_c_356_n Z Vss PM_G4_XOR2_N3_Z
cc_1 N_VSS_XI18.X0_PGD N_VDD_XI20.X0_PGD 3.18967e-19
cc_2 N_VSS_XI22.X0_PGD N_VDD_XI20.X0_PGD 0.00194647f
cc_3 N_VSS_XI18.X0_PGD N_VDD_XI16.X0_PGD 0.00196596f
cc_4 N_VSS_c_4_p N_VDD_c_96_n 0.00194647f
cc_5 N_VSS_c_5_p N_VDD_c_97_n 0.00196596f
cc_6 N_VSS_c_6_p N_VDD_c_98_n 3.76525e-19
cc_7 N_VSS_c_7_p N_VDD_c_99_n 9.5668e-19
cc_8 N_VSS_c_8_p N_VDD_c_99_n 0.00165395f
cc_9 N_VSS_c_9_p N_VDD_c_99_n 0.00452338f
cc_10 N_VSS_c_10_p N_VDD_c_99_n 0.00889981f
cc_11 N_VSS_c_11_p N_VDD_c_99_n 9.16632e-19
cc_12 N_VSS_XI18.X0_PGD N_VDD_c_104_n 3.80615e-19
cc_13 N_VSS_c_13_p N_VDD_c_104_n 4.35319e-19
cc_14 N_VSS_c_14_p N_VDD_c_104_n 3.66936e-19
cc_15 N_VSS_c_10_p N_VDD_c_104_n 0.0039632f
cc_16 N_VSS_c_7_p N_VDD_c_108_n 2.57623e-19
cc_17 N_VSS_c_8_p N_VDD_c_108_n 3.02798e-19
cc_18 N_VSS_c_18_p N_VDD_c_108_n 0.00357068f
cc_19 N_VSS_c_19_p N_VDD_c_111_n 0.00106367f
cc_20 N_VSS_c_8_p N_VDD_c_112_n 4.43088e-19
cc_21 N_VSS_c_5_p N_VDD_c_113_n 3.89167e-19
cc_22 N_VSS_c_22_p N_VDD_c_113_n 3.89167e-19
cc_23 N_VSS_c_13_p N_VDD_c_113_n 0.00161703f
cc_24 N_VSS_c_14_p N_VDD_c_113_n 2.26455e-19
cc_25 N_VSS_c_25_p N_VDD_c_113_n 0.00348402f
cc_26 N_VSS_c_26_p N_VDD_c_113_n 0.00600907f
cc_27 N_VSS_c_27_p N_VDD_c_113_n 7.74609e-19
cc_28 N_VSS_c_28_p N_VDD_c_120_n 0.00107963f
cc_29 N_VSS_c_29_p N_VDD_c_121_n 9.20609e-19
cc_30 N_VSS_c_30_p N_VDD_c_121_n 3.82294e-19
cc_31 N_VSS_c_4_p N_VDD_c_123_n 3.76472e-19
cc_32 N_VSS_c_29_p N_VDD_c_123_n 0.00141228f
cc_33 N_VSS_c_30_p N_VDD_c_123_n 0.00112249f
cc_34 N_VSS_c_18_p N_VDD_c_123_n 0.00616046f
cc_35 N_VSS_c_13_p N_VDD_c_127_n 9.25616e-19
cc_36 N_VSS_c_36_p N_VDD_c_127_n 8.475e-19
cc_37 N_VSS_c_14_p N_VDD_c_127_n 3.99794e-19
cc_38 N_VSS_c_38_p N_VDD_c_130_n 2.88732e-19
cc_39 N_VSS_c_29_p N_VDD_c_130_n 0.00232715f
cc_40 N_VSS_c_30_p N_VDD_c_130_n 9.55109e-19
cc_41 N_VSS_c_41_p N_VDD_c_133_n 9.21122e-19
cc_42 N_VSS_c_10_p N_VDD_c_134_n 0.0010705f
cc_43 N_VSS_c_18_p N_VDD_c_135_n 9.68246e-19
cc_44 N_VSS_c_29_p N_VDD_c_136_n 3.48267e-19
cc_45 N_VSS_c_30_p N_VDD_c_136_n 8.00903e-19
cc_46 N_VSS_c_13_p N_VDD_c_138_n 3.48267e-19
cc_47 N_VSS_c_14_p N_VDD_c_138_n 6.489e-19
cc_48 N_VSS_XI18.X0_PGD N_A_c_191_n 4.09718e-19
cc_49 N_VSS_XI22.X0_PGD N_A_c_191_n 2.49973e-19
cc_50 N_VSS_c_14_p N_A_c_193_n 5.35095e-19
cc_51 N_VSS_XI22.X0_PGD N_A_c_194_n 2.49973e-19
cc_52 N_VSS_c_14_p N_A_c_195_n 2.15082e-19
cc_53 N_VSS_c_36_p N_A_c_196_n 0.00705874f
cc_54 N_VSS_c_10_p N_A_c_196_n 9.14669e-19
cc_55 N_VSS_c_55_p N_A_c_196_n 0.00173435f
cc_56 N_VSS_c_41_p N_A_c_196_n 3.96468e-19
cc_57 N_VSS_c_57_p N_A_c_196_n 4.40676e-19
cc_58 N_VSS_c_55_p N_A_c_201_n 6.19395e-19
cc_59 N_VSS_c_13_p N_A_c_202_n 2.15082e-19
cc_60 N_VSS_c_55_p N_A_c_203_n 4.24683e-19
cc_61 N_VSS_c_7_p N_NET1_c_245_n 3.43419e-19
cc_62 N_VSS_c_8_p N_NET1_c_246_n 0.00115894f
cc_63 N_VSS_c_29_p N_NET1_c_247_n 0.00149535f
cc_64 N_VSS_c_9_p N_NET1_c_248_n 7.76947e-19
cc_65 N_VSS_c_18_p N_NET1_c_248_n 6.52479e-19
cc_66 N_VSS_c_6_p N_NET2_c_279_n 3.43419e-19
cc_67 N_VSS_c_36_p N_NET2_c_279_n 3.48267e-19
cc_68 N_VSS_c_6_p N_NET2_c_281_n 3.48267e-19
cc_69 N_VSS_c_36_p N_NET2_c_281_n 0.00192385f
cc_70 N_VSS_c_10_p N_NET2_c_281_n 8.02212e-19
cc_71 N_VSS_c_36_p N_NET2_c_284_n 0.00186158f
cc_72 N_VSS_c_26_p N_NET2_c_284_n 0.00117864f
cc_73 N_VSS_c_55_p N_NET2_c_284_n 0.00504587f
cc_74 N_VSS_c_57_p N_NET2_c_284_n 0.00115623f
cc_75 N_VSS_c_13_p N_NET2_c_288_n 5.67902e-19
cc_76 N_VSS_c_26_p N_NET2_c_288_n 4.84133e-19
cc_77 N_VSS_c_30_p N_B_XI22.X0_CG 0.00322194f
cc_78 N_VSS_XI22.X0_PGD N_B_XI21.X0_PGD 0.00189584f
cc_79 N_VSS_XI18.X0_PGD N_B_c_323_n 2.60477e-19
cc_80 N_VSS_XI22.X0_PGD N_B_c_323_n 4.09718e-19
cc_81 N_VSS_XI22.X0_PGD N_B_c_325_n 4.09718e-19
cc_82 N_VSS_c_30_p N_B_c_326_n 2.76939e-19
cc_83 N_VSS_c_38_p N_B_c_327_n 0.00167898f
cc_84 N_VSS_c_6_p N_Z_c_352_n 3.43419e-19
cc_85 N_VSS_c_85_p N_Z_c_352_n 3.43419e-19
cc_86 N_VSS_c_36_p N_Z_c_352_n 3.48267e-19
cc_87 N_VSS_c_87_p N_Z_c_352_n 3.48267e-19
cc_88 N_VSS_c_6_p N_Z_c_356_n 3.48267e-19
cc_89 N_VSS_c_85_p N_Z_c_356_n 3.48267e-19
cc_90 N_VSS_c_36_p N_Z_c_356_n 4.84964e-19
cc_91 N_VSS_c_87_p N_Z_c_356_n 5.71987e-19
cc_92 N_VSS_c_55_p N_Z_c_356_n 3.20264e-19
cc_93 N_VDD_XI16.X0_PGD N_A_XI19.X0_PGD 0.00169921f
cc_94 N_VDD_XI20.X0_PGD N_A_c_191_n 2.49973e-19
cc_95 N_VDD_XI16.X0_PGD N_A_c_191_n 4.09718e-19
cc_96 N_VDD_XI16.X0_PGD N_A_c_194_n 4.09718e-19
cc_97 N_VDD_c_144_p N_A_c_208_n 0.00169921f
cc_98 N_VDD_c_99_n N_A_c_195_n 5.04211e-19
cc_99 N_VDD_c_127_n N_A_c_196_n 5.50187e-19
cc_100 N_VDD_c_138_n N_A_c_196_n 3.5189e-19
cc_101 N_VDD_c_148_p N_A_c_201_n 5.4427e-19
cc_102 N_VDD_c_99_n N_A_c_202_n 6.25289e-19
cc_103 N_VDD_c_136_n N_A_c_202_n 2.53697e-19
cc_104 N_VDD_c_127_n N_A_c_215_n 4.08069e-19
cc_105 N_VDD_c_138_n N_A_c_215_n 6.61916e-19
cc_106 N_VDD_c_148_p N_A_c_203_n 7.25922e-19
cc_107 N_VDD_c_148_p N_NET1_c_250_n 8.20153e-19
cc_108 N_VDD_c_155_p N_NET1_c_250_n 4.09731e-19
cc_109 N_VDD_c_98_n N_NET1_c_245_n 3.43419e-19
cc_110 N_VDD_c_98_n N_NET1_c_246_n 3.48267e-19
cc_111 N_VDD_c_123_n N_NET1_c_246_n 2.9283e-19
cc_112 N_VDD_c_130_n N_NET1_c_246_n 0.00152282f
cc_113 N_VDD_c_130_n N_NET1_c_247_n 0.00160739f
cc_114 N_VDD_c_148_p N_NET1_c_247_n 0.00374811f
cc_115 N_VDD_c_155_p N_NET1_c_247_n 8.18723e-19
cc_116 N_VDD_c_130_n N_NET1_c_259_n 2.78343e-19
cc_117 N_VDD_c_148_p N_NET1_c_259_n 2.37583e-19
cc_118 N_VDD_c_155_p N_NET1_c_259_n 3.70842e-19
cc_119 N_VDD_c_121_n N_NET1_c_248_n 2.88872e-19
cc_120 N_VDD_c_167_p N_NET2_c_279_n 3.67949e-19
cc_121 N_VDD_c_112_n N_NET2_c_279_n 3.72199e-19
cc_122 N_VDD_c_167_p N_NET2_c_281_n 3.9802e-19
cc_123 N_VDD_c_112_n N_NET2_c_281_n 5.226e-19
cc_124 N_VDD_c_113_n N_NET2_c_281_n 3.21336e-19
cc_125 N_VDD_c_127_n N_NET2_c_284_n 3.20822e-19
cc_126 N_VDD_c_99_n N_B_XI20.X0_CG 3.86879e-19
cc_127 N_VDD_c_136_n N_B_XI20.X0_CG 0.00180351f
cc_128 N_VDD_XI20.X0_PGD N_B_c_323_n 4.09718e-19
cc_129 N_VDD_XI16.X0_PGD N_B_c_323_n 2.60477e-19
cc_130 N_VDD_XI16.X0_PGD N_B_c_325_n 2.60477e-19
cc_131 N_VDD_c_130_n N_B_c_327_n 3.02511e-19
cc_132 N_VDD_c_148_p N_B_c_327_n 9.69761e-19
cc_133 N_VDD_c_138_n N_B_c_335_n 4.47793e-19
cc_134 N_VDD_c_98_n N_Z_c_361_n 3.43419e-19
cc_135 N_VDD_c_130_n N_Z_c_361_n 3.48267e-19
cc_136 N_VDD_c_148_p N_Z_c_361_n 2.57623e-19
cc_137 N_VDD_c_133_n N_Z_c_361_n 3.72199e-19
cc_138 N_VDD_c_185_p N_Z_c_361_n 3.43419e-19
cc_139 N_VDD_c_98_n N_Z_c_356_n 3.48267e-19
cc_140 N_VDD_c_130_n N_Z_c_356_n 7.9714e-19
cc_141 N_VDD_c_148_p N_Z_c_356_n 4.72042e-19
cc_142 N_VDD_c_133_n N_Z_c_356_n 8.30519e-19
cc_143 N_VDD_c_185_p N_Z_c_356_n 3.48267e-19
cc_144 N_A_XI23.X0_CG N_NET1_XI23.X0_PGD 9.16948e-19
cc_145 N_A_c_219_p N_NET1_XI23.X0_PGD 9.43732e-19
cc_146 N_A_c_201_n N_NET1_c_247_n 0.00175052f
cc_147 N_A_c_203_n N_NET1_c_247_n 5.83558e-19
cc_148 N_A_XI23.X0_CG N_NET1_c_259_n 0.00320789f
cc_149 N_A_c_219_p N_NET1_c_259_n 4.20251e-19
cc_150 N_A_XI23.X0_CG N_NET2_XI21.X0_CG 2.29068e-19
cc_151 N_A_XI19.X0_PGD N_NET2_XI17.X0_PGD 0.00174694f
cc_152 N_A_c_194_n N_NET2_XI17.X0_PGD 3.14428e-19
cc_153 N_A_c_219_p N_NET2_XI17.X0_PGD 3.71891e-19
cc_154 N_A_XI19.X0_PGD N_NET2_c_300_n 4.64512e-19
cc_155 N_A_c_208_n N_NET2_c_301_n 0.00174694f
cc_156 N_A_c_191_n N_NET2_c_279_n 6.03094e-19
cc_157 N_A_c_196_n N_NET2_c_284_n 0.002281f
cc_158 N_A_c_201_n N_NET2_c_284_n 9.32615e-19
cc_159 N_A_c_215_n N_NET2_c_284_n 3.44698e-19
cc_160 N_A_c_196_n N_NET2_c_306_n 3.44698e-19
cc_161 N_A_c_215_n N_NET2_c_306_n 6.78604e-19
cc_162 N_A_c_194_n N_B_XI19.X0_CG 0.003858f
cc_163 N_A_c_191_n N_B_c_323_n 0.00635057f
cc_164 N_A_c_202_n N_B_c_338_n 9.89912e-19
cc_165 N_A_c_194_n N_B_c_325_n 0.00470625f
cc_166 N_A_c_194_n N_B_c_340_n 0.00225174f
cc_167 N_A_c_191_n N_B_c_335_n 0.00106939f
cc_168 N_A_c_196_n N_Z_c_356_n 0.00384185f
cc_169 N_A_c_201_n N_Z_c_356_n 0.00366674f
cc_170 N_A_c_219_p N_Z_c_356_n 9.50702e-19
cc_171 N_NET1_XI23.X0_PGD N_NET2_XI21.X0_CG 2.3921e-19
cc_172 N_NET1_c_270_p N_NET2_XI17.X0_PGD 0.00794356f
cc_173 N_NET1_XI23.X0_PGD N_NET2_c_300_n 0.00388625f
cc_174 N_NET1_c_245_n N_NET2_c_279_n 2.80316e-19
cc_175 N_NET1_XI23.X0_PGD N_B_XI21.X0_PGD 0.00215617f
cc_176 N_NET1_XI17.X0_CG N_B_XI19.X0_CG 2.58346e-19
cc_177 N_NET1_c_245_n N_B_c_323_n 5.56563e-19
cc_178 N_NET1_c_270_p N_B_c_340_n 2.58346e-19
cc_179 N_NET1_c_250_n N_B_c_327_n 0.00193019f
cc_180 N_NET1_c_247_n N_Z_c_356_n 2.27374e-19
cc_181 N_NET2_XI21.X0_CG N_B_XI21.X0_PGD 0.00204226f
cc_182 N_NET2_c_300_n N_B_XI21.X0_PGD 0.00163867f
cc_183 N_NET2_XI17.X0_PGD N_B_c_340_n 0.00351134f
cc_184 N_NET2_c_315_p N_B_c_340_n 0.00405072f
cc_185 N_NET2_c_300_n N_Z_c_361_n 7.50005e-19
cc_186 N_NET2_c_300_n N_Z_c_352_n 2.48148e-19
cc_187 N_NET2_XI17.X0_PGD N_Z_c_356_n 0.00113722f
cc_188 N_NET2_c_300_n N_Z_c_356_n 2.5304e-19
cc_189 N_NET2_c_284_n N_Z_c_356_n 3.45637e-19
cc_190 N_B_c_340_n N_Z_c_356_n 0.00106974f
*
.ends
*
*
.subckt XOR2_HPNW12 A B Y VDD VSS
xgate (VSS VDD A B Y) G4_XOR2_N3
.ends
*
* File: G5_XOR3_N3.pex.netlist
* Created: Fri Apr  1 15:48:12 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XOR3_N3_VDD 2 5 9 12 14 17 34 35 44 45 54 55 65 69 74 77 79 80 81
+ 84 86 90 93 96 98 102 104 108 112 114 116 118 119 125 134 139 Vss
c113 139 Vss 0.00510833f
c114 134 Vss 0.00495479f
c115 125 Vss 0.00566756f
c116 119 Vss 2.39889e-19
c117 118 Vss 4.92173e-19
c118 117 Vss 5.50975e-19
c119 114 Vss 4.52364e-19
c120 112 Vss 0.00180866f
c121 108 Vss 0.00116218f
c122 104 Vss 0.00632073f
c123 102 Vss 0.0010418f
c124 98 Vss 0.00598007f
c125 96 Vss 0.00126332f
c126 93 Vss 0.00323042f
c127 90 Vss 0.00584753f
c128 86 Vss 0.00654417f
c129 84 Vss 0.00154142f
c130 81 Vss 8.68392e-19
c131 80 Vss 0.00938293f
c132 79 Vss 0.0122224f
c133 77 Vss 0.00304889f
c134 74 Vss 0.00820121f
c135 69 Vss 0.00836757f
c136 65 Vss 0.00811483f
c137 55 Vss 0.0356247f
c138 54 Vss 0.10084f
c139 45 Vss 0.0356281f
c140 44 Vss 0.101312f
c141 35 Vss 0.0346562f
c142 34 Vss 0.0991017f
c143 17 Vss 0.378774f
c144 9 Vss 0.379342f
c145 5 Vss 0.383323f
r146 110 112 6.16843
r147 108 139 1.16709
r148 106 108 2.16729
r149 105 119 0.494161
r150 104 110 0.652036
r151 104 105 7.46046
r152 102 134 1.16709
r153 100 119 0.128424
r154 100 102 2.16729
r155 99 118 0.494161
r156 98 106 0.652036
r157 98 99 10.3363
r158 94 117 0.0828784
r159 94 96 2.00578
r160 93 118 0.128424
r161 92 117 0.551426
r162 92 93 5.50157
r163 90 125 1.16709
r164 88 117 0.551426
r165 88 90 7.66886
r166 87 116 0.326018
r167 86 118 0.494161
r168 86 87 10.1279
r169 82 114 0.0828784
r170 82 84 1.82344
r171 80 119 0.494161
r172 80 81 15.8795
r173 79 116 0.326018
r174 78 114 0.551426
r175 78 79 18.3386
r176 77 114 0.551426
r177 76 81 0.652036
r178 76 77 5.50157
r179 74 112 1.16709
r180 69 96 1.16709
r181 65 84 1.16709
r182 57 139 0.0476429
r183 55 57 1.45875
r184 54 58 0.652036
r185 54 57 1.45875
r186 51 55 0.652036
r187 47 134 0.0476429
r188 45 47 1.45875
r189 44 48 0.652036
r190 44 47 1.45875
r191 41 45 0.652036
r192 37 125 0.238214
r193 35 37 1.45875
r194 34 38 0.652036
r195 34 37 1.45875
r196 31 35 0.652036
r197 17 58 5.1348
r198 17 51 5.1348
r199 14 74 0.123773
r200 12 69 0.123773
r201 9 48 5.1348
r202 9 41 5.1348
r203 5 38 5.1348
r204 5 31 5.1348
r205 2 65 0.123773
.ends

.subckt PM_G5_XOR3_N3_C 2 4 6 8 17 20 23 32 37 40 44 47 52 57 84 92 98 Vss
c49 98 Vss 3.22849e-19
c50 92 Vss 0.00543331f
c51 84 Vss 0.00847968f
c52 57 Vss 0.004971f
c53 52 Vss 7.31044e-19
c54 47 Vss 9.97921e-19
c55 40 Vss 0.00163759f
c56 37 Vss 0.0082356f
c57 32 Vss 0.00958317f
c58 23 Vss 2.04877e-19
c59 20 Vss 0.221837f
c60 17 Vss 0.180502f
c61 15 Vss 0.0247918f
c62 4 Vss 0.188411f
r63 93 98 0.441572
r64 92 94 0.655813
r65 92 93 9.04425
r66 88 98 0.174814
r67 84 98 0.441572
r68 52 94 3.33429
r69 47 88 3.33429
r70 40 57 1.16709
r71 40 84 22.1365
r72 40 44 0.0416786
r73 37 52 1.16709
r74 32 47 1.16709
r75 23 57 0.0476429
r76 21 23 0.326018
r77 21 23 0.1167
r78 20 24 0.652036
r79 20 23 6.7686
r80 17 57 0.357321
r81 15 23 0.326018
r82 15 17 0.40845
r83 8 37 0.123773
r84 6 32 0.123773
r85 4 24 5.1348
r86 2 17 4.72635
.ends

.subckt PM_G5_XOR3_N3_VSS 3 6 8 11 15 18 34 37 44 45 54 55 57 66 70 73 78 83 88
+ 93 98 107 112 121 123 124 125 130 131 136 142 145 154 155 156 Vss
c110 156 Vss 3.75522e-19
c111 155 Vss 3.91906e-19
c112 154 Vss 4.4306e-19
c113 142 Vss 0.00252991f
c114 136 Vss 0.00380695f
c115 131 Vss 8.45126e-19
c116 130 Vss 0.00638861f
c117 125 Vss 8.42189e-19
c118 124 Vss 0.0059194f
c119 123 Vss 0.00432257f
c120 121 Vss 0.00374747f
c121 112 Vss 0.00407665f
c122 107 Vss 0.00420294f
c123 98 Vss 0.00605485f
c124 93 Vss 0.00198064f
c125 88 Vss 8.56162e-19
c126 83 Vss 0.00102135f
c127 78 Vss 0.00266782f
c128 73 Vss 0.00352975f
c129 70 Vss 0.0100681f
c130 66 Vss 0.00715185f
c131 57 Vss 9.01088e-20
c132 55 Vss 0.0347733f
c133 54 Vss 0.0999406f
c134 45 Vss 0.035088f
c135 44 Vss 0.0994129f
c136 37 Vss 5.39995e-20
c137 35 Vss 0.0349058f
c138 34 Vss 0.100344f
c139 15 Vss 0.379408f
c140 11 Vss 0.379783f
c141 8 Vss 0.00143493f
c142 3 Vss 0.3841f
r143 143 156 0.494161
r144 143 145 6.62689
r145 142 150 0.652036
r146 142 145 0.833571
r147 138 156 0.128424
r148 137 155 0.494161
r149 136 146 0.652036
r150 136 137 7.46046
r151 132 155 0.128424
r152 130 156 0.494161
r153 130 131 15.8795
r154 126 154 0.0828784
r155 124 155 0.494161
r156 124 125 13.0037
r157 123 131 0.652036
r158 122 154 0.551426
r159 122 123 13.8373
r160 121 154 0.551426
r161 120 125 0.652036
r162 120 121 10.0029
r163 93 150 6.16843
r164 88 112 1.16709
r165 88 146 2.16729
r166 83 107 1.16709
r167 83 138 2.16729
r168 78 132 6.16843
r169 73 98 1.16709
r170 73 126 4.33978
r171 70 93 1.16709
r172 66 78 1.16709
r173 57 112 0.0476429
r174 55 57 1.45875
r175 54 58 0.652036
r176 54 57 1.45875
r177 51 55 0.652036
r178 47 107 0.0476429
r179 45 47 1.45875
r180 44 48 0.652036
r181 44 47 1.45875
r182 41 45 0.652036
r183 37 98 0.238214
r184 35 37 1.45875
r185 34 38 0.652036
r186 34 37 1.45875
r187 31 35 0.652036
r188 18 70 0.123773
r189 15 58 5.1348
r190 15 51 5.1348
r191 11 48 5.1348
r192 11 41 5.1348
r193 8 66 0.123773
r194 6 66 0.123773
r195 3 38 5.1348
r196 3 31 5.1348
.ends

.subckt PM_G5_XOR3_N3_CI 2 4 6 8 23 26 31 34 39 44 79 80 82 84 89 Vss
c52 95 Vss 8.92453e-20
c53 89 Vss 0.00607467f
c54 84 Vss 1.6915e-19
c55 83 Vss 1.82188e-19
c56 82 Vss 0.00167496f
c57 80 Vss 4.34795e-19
c58 79 Vss 0.00544906f
c59 44 Vss 7.72828e-19
c60 39 Vss 9.91594e-19
c61 34 Vss 0.00323815f
c62 31 Vss 0.00967911f
c63 26 Vss 0.00811165f
c64 23 Vss 0.00522928f
c65 4 Vss 0.00143493f
r66 90 95 0.494161
r67 89 91 0.652036
r68 89 90 10.3363
r69 85 95 0.128424
r70 83 95 0.494161
r71 83 84 1.50043
r72 82 84 0.652036
r73 81 82 6.46018
r74 79 81 0.652036
r75 79 80 19.1721
r76 75 80 0.652036
r77 44 91 3.41764
r78 39 85 3.41764
r79 34 75 8.62746
r80 31 44 1.16709
r81 26 39 1.16709
r82 23 34 1.16709
r83 8 31 0.123773
r84 6 26 0.123773
r85 4 23 0.123773
r86 2 23 0.123773
.ends

.subckt PM_G5_XOR3_N3_A 2 4 7 11 24 44 45 49 51 54 55 57 59 62 67 72 Vss
c67 72 Vss 0.00561856f
c68 67 Vss 0.00509443f
c69 59 Vss 9.40202e-19
c70 57 Vss 0.00665603f
c71 55 Vss 6.2663e-19
c72 54 Vss 0.00565582f
c73 51 Vss 0.00800572f
c74 49 Vss 0.135088f
c75 45 Vss 0.128114f
c76 44 Vss 1.14131e-19
c77 24 Vss 0.221923f
c78 21 Vss 0.18375f
c79 19 Vss 0.0247918f
c80 7 Vss 1.43819f
c81 4 Vss 0.194116f
r82 64 67 1.16709
r83 62 64 0.0416786
r84 59 62 0.833571
r85 57 72 1.16709
r86 55 57 9.66422
r87 53 55 0.655813
r88 53 54 10.4613
r89 52 59 0.0685365
r90 51 54 0.652036
r91 51 52 10.2113
r92 47 49 4.53833
r93 44 72 0.0238214
r94 44 45 2.26917
r95 41 44 2.26917
r96 36 49 0.00605528
r97 35 45 0.00605528
r98 32 47 0.00605528
r99 31 41 0.00605528
r100 27 67 0.0952857
r101 25 27 0.326018
r102 25 27 0.1167
r103 24 28 0.652036
r104 24 27 6.7686
r105 21 27 0.3335
r106 19 27 0.326018
r107 19 21 0.2334
r108 11 36 5.1348
r109 11 32 5.1348
r110 7 11 17.9718
r111 7 35 5.1348
r112 7 11 17.9718
r113 7 31 5.1348
r114 4 28 5.1348
r115 2 21 4.9014
.ends

.subckt PM_G5_XOR3_N3_BI 2 4 6 8 18 21 29 32 37 42 51 56 65 71 72 80 Vss
c62 80 Vss 3.85169e-19
c63 72 Vss 3.10144e-19
c64 71 Vss 7.91966e-19
c65 65 Vss 0.00115548f
c66 56 Vss 0.00255458f
c67 51 Vss 0.0023957f
c68 42 Vss 0.00128972f
c69 37 Vss 0.00247226f
c70 32 Vss 0.00178645f
c71 29 Vss 0.00520864f
c72 21 Vss 0.166484f
c73 6 Vss 0.166668f
c74 4 Vss 0.00143493f
r75 76 80 0.655813
r76 71 72 0.655813
r77 70 71 3.501
r78 65 70 0.655813
r79 42 56 1.16709
r80 42 72 2.00578
r81 37 51 1.16709
r82 37 80 12.0712
r83 37 65 2.00578
r84 32 76 3.33429
r85 29 32 1.16709
r86 21 56 0.50025
r87 18 51 0.50025
r88 8 21 4.37625
r89 6 18 4.37625
r90 4 29 0.123773
r91 2 29 0.123773
.ends

.subckt PM_G5_XOR3_N3_AI 2 4 7 11 31 37 43 46 51 60 73 79 Vss
c44 79 Vss 2.91008e-19
c45 73 Vss 0.00515518f
c46 60 Vss 0.0064096f
c47 51 Vss 0.00263851f
c48 46 Vss 0.0021137f
c49 43 Vss 0.0046119f
c50 37 Vss 0.12791f
c51 31 Vss 0.131715f
c52 7 Vss 1.42572f
c53 4 Vss 0.00143493f
r54 75 79 0.652036
r55 73 79 13.7539
r56 51 60 1.16709
r57 51 73 2.75079
r58 46 75 6.16843
r59 43 46 1.16709
r60 36 60 0.0238214
r61 36 37 2.334
r62 33 36 2.20433
r63 29 31 4.53833
r64 26 37 0.00605528
r65 25 31 0.00605528
r66 22 33 0.00605528
r67 21 29 0.00605528
r68 11 26 5.1348
r69 11 22 5.1348
r70 7 11 17.9718
r71 7 25 5.1348
r72 7 11 17.9718
r73 7 21 5.1348
r74 4 43 0.123773
r75 2 43 0.123773
.ends

.subckt PM_G5_XOR3_N3_B 2 4 6 8 16 17 24 26 33 38 42 45 50 55 60 65 73 74 80 86
+ 91 92 Vss
c69 92 Vss 2.0377e-19
c70 91 Vss 6.9543e-19
c71 86 Vss 8.47373e-19
c72 80 Vss 9.51093e-19
c73 74 Vss 5.10711e-19
c74 73 Vss 0.00481884f
c75 65 Vss 0.00266055f
c76 60 Vss 0.00231285f
c77 55 Vss 0.00437951f
c78 50 Vss 0.00146415f
c79 45 Vss 4.84439e-19
c80 42 Vss 7.72719e-19
c81 38 Vss 7.58106e-19
c82 33 Vss 9.01088e-20
c83 26 Vss 0.166484f
c84 24 Vss 1.01938e-19
c85 20 Vss 0.0247918f
c86 17 Vss 0.0340157f
c87 16 Vss 0.186033f
c88 8 Vss 0.166484f
c89 4 Vss 0.180512f
c90 2 Vss 0.191454f
r91 90 92 0.655813
r92 90 91 3.501
r93 86 91 0.655813
r94 73 80 0.0685365
r95 73 74 10.3363
r96 69 74 0.652036
r97 50 65 1.16709
r98 50 92 2.00578
r99 45 60 1.16709
r100 45 86 2.00578
r101 45 80 2.04225
r102 38 55 1.16709
r103 38 69 2.20896
r104 38 42 0.0729375
r105 36 55 0.0476429
r106 33 65 0.50025
r107 26 60 0.50025
r108 24 55 0.357321
r109 20 36 0.326018
r110 20 24 0.40845
r111 17 36 6.7686
r112 16 36 0.326018
r113 16 36 0.1167
r114 13 17 0.652036
r115 8 33 4.37625
r116 6 26 4.37625
r117 4 24 4.72635
r118 2 13 5.1348
.ends

.subckt PM_G5_XOR3_N3_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00377706f
c33 27 Vss 0.00795274f
c34 23 Vss 0.00720799f
c35 8 Vss 0.00143493f
c36 6 Vss 0.00334888f
r37 33 35 7.21039
r38 30 40 1.16709
r39 30 33 5.62661
r40 27 35 1.16709
r41 23 40 0.05
r42 8 27 0.123773
r43 6 23 0.123773
r44 4 27 0.123773
r45 2 23 0.123773
.ends

.subckt G5_XOR3_N3  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI25.X0 N_CI_XI25.X0_D N_VSS_XI25.X0_PGD N_C_XI25.X0_CG N_VSS_XI25.X0_PGD
+ N_VDD_XI25.X0_S TIGFET_HPNW12
XI22.X0 N_CI_XI22.X0_D N_VDD_XI22.X0_PGD N_C_XI22.X0_CG N_VDD_XI22.X0_PGD
+ N_VSS_XI22.X0_S TIGFET_HPNW12
XI21.X0 N_BI_XI21.X0_D N_VDD_XI21.X0_PGD N_B_XI21.X0_CG N_VDD_XI21.X0_PGD
+ N_VSS_XI21.X0_S TIGFET_HPNW12
XI23.X0 N_AI_XI23.X0_D N_VSS_XI23.X0_PGD N_A_XI23.X0_CG N_VSS_XI23.X0_PGD
+ N_VDD_XI23.X0_S TIGFET_HPNW12
XI24.X0 N_BI_XI24.X0_D N_VSS_XI24.X0_PGD N_B_XI24.X0_CG N_VSS_XI24.X0_PGD
+ N_VDD_XI24.X0_S TIGFET_HPNW12
XI20.X0 N_AI_XI20.X0_D N_VDD_XI20.X0_PGD N_A_XI20.X0_CG N_VDD_XI20.X0_PGD
+ N_VSS_XI20.X0_S TIGFET_HPNW12
XI29.X0 N_Z_XI29.X0_D N_AI_XI29.X0_PGD N_BI_XI29.X0_CG N_AI_XI29.X0_PGD
+ N_C_XI29.X0_S TIGFET_HPNW12
XI27.X0 N_Z_XI27.X0_D N_AI_XI27.X0_PGD N_B_XI27.X0_CG N_AI_XI27.X0_PGD
+ N_CI_XI27.X0_S TIGFET_HPNW12
XI28.X0 N_Z_XI28.X0_D N_A_XI28.X0_PGD N_B_XI28.X0_CG N_A_XI28.X0_PGD
+ N_C_XI28.X0_S TIGFET_HPNW12
XI26.X0 N_Z_XI26.X0_D N_A_XI26.X0_PGD N_BI_XI26.X0_CG N_A_XI26.X0_PGD
+ N_CI_XI26.X0_S TIGFET_HPNW12
*
x_PM_G5_XOR3_N3_VDD N_VDD_XI25.X0_S N_VDD_XI22.X0_PGD N_VDD_XI21.X0_PGD
+ N_VDD_XI23.X0_S N_VDD_XI24.X0_S N_VDD_XI20.X0_PGD N_VDD_c_111_p N_VDD_c_19_p
+ N_VDD_c_24_p N_VDD_c_4_p N_VDD_c_100_p N_VDD_c_20_p N_VDD_c_74_p N_VDD_c_101_p
+ N_VDD_c_6_p N_VDD_c_7_p N_VDD_c_13_p N_VDD_c_5_p N_VDD_c_61_p N_VDD_c_29_p
+ N_VDD_c_62_p N_VDD_c_30_p N_VDD_c_16_p N_VDD_c_63_p N_VDD_c_21_p N_VDD_c_10_p
+ N_VDD_c_25_p N_VDD_c_37_p N_VDD_c_11_p N_VDD_c_57_p VDD N_VDD_c_65_p
+ N_VDD_c_69_p N_VDD_c_2_p N_VDD_c_42_p N_VDD_c_38_p Vss PM_G5_XOR3_N3_VDD
x_PM_G5_XOR3_N3_C N_C_XI25.X0_CG N_C_XI22.X0_CG N_C_XI29.X0_S N_C_XI28.X0_S
+ N_C_c_130_p N_C_c_116_n N_C_c_126_p N_C_c_119_n N_C_c_157_p N_C_c_120_n C
+ N_C_c_127_p N_C_c_159_p N_C_c_122_n N_C_c_123_n N_C_c_145_p N_C_c_146_p Vss
+ PM_G5_XOR3_N3_C
x_PM_G5_XOR3_N3_VSS N_VSS_XI25.X0_PGD N_VSS_XI22.X0_S N_VSS_XI21.X0_S
+ N_VSS_XI23.X0_PGD N_VSS_XI24.X0_PGD N_VSS_XI20.X0_S N_VSS_c_170_n
+ N_VSS_c_226_n N_VSS_c_171_n N_VSS_c_173_n N_VSS_c_174_n N_VSS_c_175_n
+ N_VSS_c_269_p N_VSS_c_177_n N_VSS_c_238_p N_VSS_c_178_n N_VSS_c_183_n
+ N_VSS_c_186_n N_VSS_c_190_n N_VSS_c_194_n N_VSS_c_195_n N_VSS_c_198_n
+ N_VSS_c_202_n N_VSS_c_206_n N_VSS_c_209_n N_VSS_c_211_n N_VSS_c_212_n
+ N_VSS_c_213_n N_VSS_c_217_n N_VSS_c_218_n N_VSS_c_221_n VSS N_VSS_c_222_n
+ N_VSS_c_223_n N_VSS_c_224_n Vss PM_G5_XOR3_N3_VSS
x_PM_G5_XOR3_N3_CI N_CI_XI25.X0_D N_CI_XI22.X0_D N_CI_XI27.X0_S N_CI_XI26.X0_S
+ N_CI_c_273_n N_CI_c_286_n N_CI_c_317_p N_CI_c_275_n N_CI_c_292_n N_CI_c_319_p
+ N_CI_c_279_n N_CI_c_295_n N_CI_c_296_n N_CI_c_308_p N_CI_c_302_p Vss
+ PM_G5_XOR3_N3_CI
x_PM_G5_XOR3_N3_A N_A_XI23.X0_CG N_A_XI20.X0_CG N_A_XI28.X0_PGD N_A_XI26.X0_PGD
+ N_A_c_325_n N_A_c_374_p N_A_c_365_p N_A_c_367_p N_A_c_326_n N_A_c_332_n
+ N_A_c_333_n N_A_c_340_n N_A_c_334_n A N_A_c_335_n N_A_c_378_p Vss
+ PM_G5_XOR3_N3_A
x_PM_G5_XOR3_N3_BI N_BI_XI21.X0_D N_BI_XI24.X0_D N_BI_XI29.X0_CG N_BI_XI26.X0_CG
+ N_BI_c_412_n N_BI_c_413_n N_BI_c_392_n N_BI_c_395_n N_BI_c_399_n N_BI_c_410_n
+ N_BI_c_418_n N_BI_c_419_n N_BI_c_402_n N_BI_c_440_p N_BI_c_428_p N_BI_c_403_n
+ Vss PM_G5_XOR3_N3_BI
x_PM_G5_XOR3_N3_AI N_AI_XI23.X0_D N_AI_XI20.X0_D N_AI_XI29.X0_PGD
+ N_AI_XI27.X0_PGD N_AI_c_465_n N_AI_c_455_n N_AI_c_456_n N_AI_c_458_n
+ N_AI_c_471_n N_AI_c_492_p N_AI_c_463_n N_AI_c_473_n Vss PM_G5_XOR3_N3_AI
x_PM_G5_XOR3_N3_B N_B_XI21.X0_CG N_B_XI24.X0_CG N_B_XI27.X0_CG N_B_XI28.X0_CG
+ N_B_c_499_n N_B_c_500_n N_B_c_507_n N_B_c_557_n N_B_c_521_n N_B_c_501_n B
+ N_B_c_537_n N_B_c_512_n N_B_c_509_n N_B_c_541_n N_B_c_529_n N_B_c_502_n
+ N_B_c_514_n N_B_c_548_n N_B_c_504_n N_B_c_554_n N_B_c_505_n Vss
+ PM_G5_XOR3_N3_B
x_PM_G5_XOR3_N3_Z N_Z_XI29.X0_D N_Z_XI27.X0_D N_Z_XI28.X0_D N_Z_XI26.X0_D
+ N_Z_c_567_n N_Z_c_574_n N_Z_c_571_n Z Vss PM_G5_XOR3_N3_Z
cc_1 N_VDD_XI21.X0_PGD N_C_XI22.X0_CG 0.00111653f
cc_2 N_VDD_c_2_p N_C_XI22.X0_CG 0.00108697f
cc_3 N_VDD_XI22.X0_PGD N_C_c_116_n 4.20258e-19
cc_4 N_VDD_c_4_p N_C_c_116_n 0.00111653f
cc_5 N_VDD_c_5_p N_C_c_116_n 0.00135138f
cc_6 N_VDD_c_6_p N_C_c_119_n 3.43419e-19
cc_7 N_VDD_c_7_p N_C_c_120_n 4.76491e-19
cc_8 N_VDD_c_5_p N_C_c_120_n 0.00161703f
cc_9 N_VDD_c_5_p N_C_c_122_n 2.84771e-19
cc_10 N_VDD_c_10_p N_C_c_123_n 5.24769e-19
cc_11 N_VDD_c_11_p N_C_c_123_n 8.43519e-19
cc_12 N_VDD_XI22.X0_PGD N_VSS_XI25.X0_PGD 0.00200994f
cc_13 N_VDD_c_13_p N_VSS_XI25.X0_PGD 4.18763e-19
cc_14 N_VDD_XI21.X0_PGD N_VSS_XI23.X0_PGD 2.44446e-19
cc_15 N_VDD_XI20.X0_PGD N_VSS_XI23.X0_PGD 0.00201012f
cc_16 N_VDD_c_16_p N_VSS_XI23.X0_PGD 4.21402e-19
cc_17 N_VDD_XI21.X0_PGD N_VSS_XI24.X0_PGD 0.00200584f
cc_18 N_VDD_XI20.X0_PGD N_VSS_XI24.X0_PGD 2.31301e-19
cc_19 N_VDD_c_19_p N_VSS_c_170_n 0.00200994f
cc_20 N_VDD_c_20_p N_VSS_c_171_n 0.00201012f
cc_21 N_VDD_c_21_p N_VSS_c_171_n 3.00545e-19
cc_22 N_VDD_c_21_p N_VSS_c_173_n 3.89167e-19
cc_23 N_VDD_c_11_p N_VSS_c_174_n 2.35465e-19
cc_24 N_VDD_c_24_p N_VSS_c_175_n 0.00200584f
cc_25 N_VDD_c_25_p N_VSS_c_175_n 3.89167e-19
cc_26 N_VDD_c_5_p N_VSS_c_177_n 2.74986e-19
cc_27 N_VDD_c_13_p N_VSS_c_178_n 4.32468e-19
cc_28 N_VDD_c_5_p N_VSS_c_178_n 3.08724e-19
cc_29 N_VDD_c_29_p N_VSS_c_178_n 0.00111881f
cc_30 N_VDD_c_30_p N_VSS_c_178_n 3.98949e-19
cc_31 N_VDD_c_2_p N_VSS_c_178_n 3.48267e-19
cc_32 N_VDD_c_5_p N_VSS_c_183_n 2.9533e-19
cc_33 N_VDD_c_10_p N_VSS_c_183_n 7.43603e-19
cc_34 N_VDD_c_11_p N_VSS_c_183_n 8.20353e-19
cc_35 N_VDD_c_16_p N_VSS_c_186_n 6.74818e-19
cc_36 N_VDD_c_21_p N_VSS_c_186_n 0.00161703f
cc_37 N_VDD_c_37_p N_VSS_c_186_n 8.6926e-19
cc_38 N_VDD_c_38_p N_VSS_c_186_n 3.48267e-19
cc_39 N_VDD_c_10_p N_VSS_c_190_n 6.78479e-19
cc_40 N_VDD_c_25_p N_VSS_c_190_n 0.00161703f
cc_41 N_VDD_c_11_p N_VSS_c_190_n 0.0024227f
cc_42 N_VDD_c_42_p N_VSS_c_190_n 3.48267e-19
cc_43 N_VDD_c_37_p N_VSS_c_194_n 7.32365e-19
cc_44 N_VDD_c_13_p N_VSS_c_195_n 4.41003e-19
cc_45 N_VDD_c_30_p N_VSS_c_195_n 3.89161e-19
cc_46 N_VDD_c_2_p N_VSS_c_195_n 7.99831e-19
cc_47 N_VDD_c_16_p N_VSS_c_198_n 3.48267e-19
cc_48 N_VDD_c_21_p N_VSS_c_198_n 2.26455e-19
cc_49 N_VDD_c_37_p N_VSS_c_198_n 3.99794e-19
cc_50 N_VDD_c_38_p N_VSS_c_198_n 6.489e-19
cc_51 N_VDD_c_10_p N_VSS_c_202_n 3.82294e-19
cc_52 N_VDD_c_25_p N_VSS_c_202_n 2.26455e-19
cc_53 N_VDD_c_11_p N_VSS_c_202_n 9.55109e-19
cc_54 N_VDD_c_42_p N_VSS_c_202_n 6.46219e-19
cc_55 N_VDD_c_7_p N_VSS_c_206_n 0.00419405f
cc_56 N_VDD_c_13_p N_VSS_c_206_n 0.00330716f
cc_57 N_VDD_c_57_p N_VSS_c_206_n 0.0010705f
cc_58 N_VDD_c_13_p N_VSS_c_209_n 0.00977753f
cc_59 N_VDD_c_30_p N_VSS_c_209_n 0.00139461f
cc_60 N_VDD_c_5_p N_VSS_c_211_n 0.0097003f
cc_61 N_VDD_c_61_p N_VSS_c_212_n 0.00107633f
cc_62 N_VDD_c_62_p N_VSS_c_213_n 0.00839359f
cc_63 N_VDD_c_63_p N_VSS_c_213_n 6.54257e-19
cc_64 N_VDD_c_21_p N_VSS_c_213_n 0.00374326f
cc_65 N_VDD_c_65_p N_VSS_c_213_n 0.00149946f
cc_66 N_VDD_c_13_p N_VSS_c_217_n 0.00107845f
cc_67 N_VDD_c_5_p N_VSS_c_218_n 0.00143483f
cc_68 N_VDD_c_25_p N_VSS_c_218_n 0.00612925f
cc_69 N_VDD_c_69_p N_VSS_c_218_n 9.53204e-19
cc_70 N_VDD_c_21_p N_VSS_c_221_n 0.00550311f
cc_71 N_VDD_c_13_p N_VSS_c_222_n 0.00112682f
cc_72 N_VDD_c_5_p N_VSS_c_223_n 0.00111918f
cc_73 N_VDD_c_21_p N_VSS_c_224_n 7.74609e-19
cc_74 N_VDD_c_74_p N_CI_c_273_n 3.43419e-19
cc_75 N_VDD_c_29_p N_CI_c_273_n 3.72199e-19
cc_76 N_VDD_c_74_p N_CI_c_275_n 3.48267e-19
cc_77 N_VDD_c_5_p N_CI_c_275_n 3.21336e-19
cc_78 N_VDD_c_29_p N_CI_c_275_n 5.226e-19
cc_79 N_VDD_c_30_p N_CI_c_275_n 0.00102111f
cc_80 N_VDD_c_30_p N_CI_c_279_n 7.25102e-19
cc_81 N_VDD_c_63_p N_CI_c_279_n 7.87445e-19
cc_82 N_VDD_XI20.X0_PGD N_A_c_325_n 3.97033e-19
cc_83 N_VDD_XI20.X0_PGD N_A_c_326_n 2.7861e-19
cc_84 N_VDD_c_6_p N_A_c_326_n 2.23042e-19
cc_85 N_VDD_c_21_p N_A_c_326_n 3.21337e-19
cc_86 N_VDD_c_37_p N_A_c_326_n 2.93421e-19
cc_87 N_VDD_c_11_p N_A_c_326_n 3.31604e-19
cc_88 N_VDD_c_38_p N_A_c_326_n 2.04325e-19
cc_89 N_VDD_c_6_p N_A_c_332_n 9.18655e-19
cc_90 N_VDD_c_11_p N_A_c_333_n 0.00704792f
cc_91 N_VDD_c_30_p N_A_c_334_n 0.00104803f
cc_92 N_VDD_c_30_p N_A_c_335_n 5.71346e-19
cc_93 N_VDD_c_6_p N_BI_c_392_n 3.43419e-19
cc_94 N_VDD_c_25_p N_BI_c_392_n 2.74986e-19
cc_95 N_VDD_c_11_p N_BI_c_392_n 3.48267e-19
cc_96 N_VDD_c_6_p N_BI_c_395_n 3.48267e-19
cc_97 N_VDD_c_25_p N_BI_c_395_n 2.9533e-19
cc_98 N_VDD_c_11_p N_BI_c_395_n 4.99861e-19
cc_99 N_VDD_XI20.X0_PGD N_AI_XI29.X0_PGD 3.2392e-19
cc_100 N_VDD_c_100_p N_AI_c_455_n 3.2392e-19
cc_101 N_VDD_c_101_p N_AI_c_456_n 3.43419e-19
cc_102 N_VDD_c_63_p N_AI_c_456_n 3.73302e-19
cc_103 N_VDD_c_101_p N_AI_c_458_n 3.48267e-19
cc_104 N_VDD_c_16_p N_AI_c_458_n 3.24512e-19
cc_105 N_VDD_c_63_p N_AI_c_458_n 5.23123e-19
cc_106 N_VDD_c_21_p N_AI_c_458_n 3.21336e-19
cc_107 N_VDD_c_37_p N_AI_c_458_n 5.55696e-19
cc_108 N_VDD_c_21_p N_AI_c_463_n 4.73141e-19
cc_109 N_VDD_XI22.X0_PGD N_B_XI21.X0_CG 0.00111821f
cc_110 N_VDD_XI21.X0_PGD N_B_c_499_n 4.01531e-19
cc_111 N_VDD_c_111_p N_B_c_500_n 0.00111821f
cc_112 N_VDD_c_30_p N_B_c_501_n 7.28643e-19
cc_113 N_VDD_c_11_p N_B_c_502_n 2.93412e-19
cc_114 N_C_c_116_n N_VSS_XI25.X0_PGD 4.20258e-19
cc_115 N_C_c_126_p N_VSS_c_226_n 2.76939e-19
cc_116 N_C_c_127_p N_VSS_c_183_n 7.31268e-19
cc_117 N_C_c_123_n N_VSS_c_183_n 0.00201674f
cc_118 N_C_c_123_n N_VSS_c_190_n 0.00162673f
cc_119 N_C_c_130_p N_VSS_c_195_n 0.0041528f
cc_120 N_C_c_120_n N_VSS_c_206_n 4.01014e-19
cc_121 N_C_c_123_n N_VSS_c_206_n 2.67373e-19
cc_122 N_C_c_120_n N_VSS_c_211_n 0.00171716f
cc_123 N_C_c_123_n N_VSS_c_211_n 0.00318423f
cc_124 N_C_c_123_n N_VSS_c_218_n 0.00194657f
cc_125 N_C_c_116_n N_CI_c_273_n 7.69306e-19
cc_126 N_C_c_123_n N_CI_c_275_n 7.41148e-19
cc_127 N_C_c_123_n N_CI_c_279_n 0.00247018f
cc_128 N_C_c_123_n N_A_c_326_n 2.96232e-19
cc_129 N_C_c_119_n N_A_c_332_n 8.20481e-19
cc_130 N_C_c_127_p N_A_c_332_n 0.00202163f
cc_131 N_C_c_123_n N_A_c_333_n 5.81147e-19
cc_132 N_C_c_127_p N_A_c_340_n 0.00128177f
cc_133 N_C_c_123_n N_A_c_340_n 4.89987e-19
cc_134 N_C_c_145_p N_A_c_340_n 0.00290875f
cc_135 N_C_c_146_p N_A_c_340_n 3.99251e-19
cc_136 N_C_c_123_n N_BI_c_395_n 7.95957e-19
cc_137 N_C_c_127_p N_BI_c_399_n 8.44326e-19
cc_138 N_C_c_123_n N_BI_c_399_n 0.00305118f
cc_139 N_C_c_145_p N_BI_c_399_n 4.85495e-19
cc_140 N_C_c_145_p N_BI_c_402_n 7.42134e-19
cc_141 N_C_c_123_n N_BI_c_403_n 5.13569e-19
cc_142 N_C_c_127_p N_B_c_502_n 6.36664e-19
cc_143 N_C_c_145_p N_B_c_504_n 3.34841e-19
cc_144 N_C_c_145_p N_B_c_505_n 0.0012842f
cc_145 N_C_c_119_n N_Z_c_567_n 3.43419e-19
cc_146 N_C_c_157_p N_Z_c_567_n 3.43419e-19
cc_147 N_C_c_127_p N_Z_c_567_n 3.48267e-19
cc_148 N_C_c_159_p N_Z_c_567_n 3.48267e-19
cc_149 N_C_c_157_p N_Z_c_571_n 3.48267e-19
cc_150 N_C_c_127_p N_Z_c_571_n 6.09821e-19
cc_151 N_C_c_159_p N_Z_c_571_n 5.71987e-19
cc_152 N_VSS_c_177_n N_CI_c_273_n 3.43419e-19
cc_153 N_VSS_c_183_n N_CI_c_273_n 3.48267e-19
cc_154 N_VSS_c_238_p N_CI_c_286_n 3.43419e-19
cc_155 N_VSS_c_177_n N_CI_c_275_n 3.48267e-19
cc_156 N_VSS_c_178_n N_CI_c_275_n 5.88914e-19
cc_157 N_VSS_c_183_n N_CI_c_275_n 8.10527e-19
cc_158 N_VSS_c_206_n N_CI_c_275_n 7.39772e-19
cc_159 N_VSS_c_209_n N_CI_c_275_n 9.66332e-19
cc_160 N_VSS_c_194_n N_CI_c_292_n 8.792e-19
cc_161 N_VSS_c_186_n N_CI_c_279_n 3.71583e-19
cc_162 N_VSS_c_221_n N_CI_c_279_n 4.92938e-19
cc_163 N_VSS_c_213_n N_CI_c_295_n 0.00161605f
cc_164 N_VSS_c_194_n N_CI_c_296_n 0.00179737f
cc_165 N_VSS_XI23.X0_PGD N_A_c_325_n 3.97033e-19
cc_166 N_VSS_c_194_n N_A_c_326_n 6.39942e-19
cc_167 N_VSS_c_221_n N_A_c_326_n 3.79499e-19
cc_168 N_VSS_c_198_n N_A_c_334_n 2.09367e-19
cc_169 N_VSS_c_186_n N_A_c_335_n 2.04211e-19
cc_170 N_VSS_c_198_n N_A_c_335_n 4.89964e-19
cc_171 N_VSS_c_177_n N_BI_c_392_n 3.43419e-19
cc_172 N_VSS_c_177_n N_BI_c_395_n 3.48267e-19
cc_173 N_VSS_c_183_n N_BI_c_395_n 8.48361e-19
cc_174 N_VSS_XI24.X0_PGD N_AI_XI29.X0_PGD 2.79882e-19
cc_175 N_VSS_c_174_n N_AI_c_465_n 2.79882e-19
cc_176 N_VSS_c_238_p N_AI_c_456_n 3.43419e-19
cc_177 N_VSS_c_238_p N_AI_c_458_n 3.48267e-19
cc_178 N_VSS_c_186_n N_AI_c_458_n 0.00108072f
cc_179 N_VSS_c_194_n N_AI_c_458_n 0.00227024f
cc_180 N_VSS_c_209_n N_AI_c_458_n 7.83107e-19
cc_181 N_VSS_c_194_n N_AI_c_471_n 0.00125351f
cc_182 N_VSS_c_221_n N_AI_c_463_n 0.00560835f
cc_183 N_VSS_c_221_n N_AI_c_473_n 0.00192498f
cc_184 N_VSS_XI24.X0_PGD N_B_c_499_n 4.01531e-19
cc_185 N_VSS_c_269_p N_B_c_507_n 5.35095e-19
cc_186 N_VSS_c_202_n B 2.15082e-19
cc_187 N_VSS_c_190_n N_B_c_509_n 2.15082e-19
cc_188 N_VSS_c_194_n N_B_c_502_n 2.6453e-19
cc_189 N_CI_c_279_n N_A_c_326_n 0.00190043f
cc_190 N_CI_c_279_n N_A_c_334_n 3.93937e-19
cc_191 N_CI_c_275_n N_BI_c_395_n 0.00116552f
cc_192 N_CI_c_292_n N_BI_c_399_n 2.45753e-19
cc_193 N_CI_c_279_n N_BI_c_399_n 0.00333331f
cc_194 N_CI_c_302_p N_BI_c_410_n 7.0273e-19
cc_195 N_CI_c_279_n N_BI_c_403_n 0.00154189f
cc_196 N_CI_c_279_n N_AI_c_458_n 9.328e-19
cc_197 N_CI_c_296_n N_AI_c_458_n 0.00145606f
cc_198 N_CI_c_302_p N_AI_c_471_n 0.00147513f
cc_199 N_CI_c_279_n N_AI_c_463_n 0.00163581f
cc_200 N_CI_c_308_p N_AI_c_463_n 0.00486757f
cc_201 N_CI_c_302_p N_AI_c_463_n 0.00259545f
cc_202 N_CI_c_275_n N_B_c_501_n 5.60809e-19
cc_203 N_CI_c_302_p N_B_c_512_n 5.08667e-19
cc_204 N_CI_c_292_n N_B_c_502_n 7.44351e-19
cc_205 N_CI_c_279_n N_B_c_514_n 0.00125143f
cc_206 N_CI_c_279_n N_B_c_504_n 4.54745e-19
cc_207 N_CI_c_302_p N_B_c_504_n 0.00126146f
cc_208 N_CI_c_286_n N_Z_c_574_n 3.43419e-19
cc_209 N_CI_c_317_p N_Z_c_574_n 3.43419e-19
cc_210 N_CI_c_292_n N_Z_c_574_n 3.48267e-19
cc_211 N_CI_c_319_p N_Z_c_574_n 3.48267e-19
cc_212 N_CI_c_286_n N_Z_c_571_n 3.48267e-19
cc_213 N_CI_c_317_p N_Z_c_571_n 3.48267e-19
cc_214 N_CI_c_292_n N_Z_c_571_n 5.71987e-19
cc_215 N_CI_c_319_p N_Z_c_571_n 5.71987e-19
cc_216 N_CI_c_279_n N_Z_c_571_n 6.3795e-19
cc_217 N_A_c_340_n N_BI_c_412_n 2.09474e-19
cc_218 N_A_XI28.X0_PGD N_BI_c_413_n 9.65637e-19
cc_219 N_A_c_326_n N_BI_c_395_n 3.45209e-19
cc_220 N_A_c_332_n N_BI_c_395_n 6.2874e-19
cc_221 N_A_c_332_n N_BI_c_399_n 0.00115936f
cc_222 N_A_c_340_n N_BI_c_399_n 6.34965e-19
cc_223 N_A_c_332_n N_BI_c_418_n 3.37713e-19
cc_224 N_A_XI28.X0_PGD N_BI_c_419_n 0.00133285f
cc_225 N_A_c_340_n N_BI_c_402_n 7.80641e-19
cc_226 N_A_c_326_n N_BI_c_403_n 4.18438e-19
cc_227 N_A_XI28.X0_PGD N_AI_XI29.X0_PGD 0.0174159f
cc_228 N_A_c_332_n N_AI_XI29.X0_PGD 9.45724e-19
cc_229 N_A_c_340_n N_AI_XI29.X0_PGD 7.67512e-19
cc_230 N_A_c_365_p N_AI_c_465_n 0.00199603f
cc_231 N_A_c_340_n N_AI_c_465_n 0.00129811f
cc_232 N_A_c_367_p N_AI_c_455_n 0.00201004f
cc_233 N_A_c_325_n N_AI_c_456_n 6.90199e-19
cc_234 N_A_c_326_n N_AI_c_458_n 5.93425e-19
cc_235 N_A_XI28.X0_PGD N_B_XI28.X0_CG 9.65637e-19
cc_236 N_A_c_325_n N_B_c_499_n 0.00358744f
cc_237 N_A_c_326_n N_B_c_499_n 8.32052e-19
cc_238 N_A_c_335_n N_B_c_500_n 7.41063e-19
cc_239 N_A_c_374_p N_B_c_521_n 5.35095e-19
cc_240 N_A_c_332_n N_B_c_501_n 6.26711e-19
cc_241 N_A_c_326_n B 8.224e-19
cc_242 N_A_c_332_n B 5.04818e-19
cc_243 N_A_c_378_p N_B_c_512_n 2.15082e-19
cc_244 N_A_c_325_n N_B_c_509_n 0.00108715f
cc_245 N_A_c_326_n N_B_c_509_n 6.90512e-19
cc_246 N_A_c_332_n N_B_c_509_n 6.85754e-19
cc_247 N_A_XI28.X0_PGD N_B_c_529_n 0.00133285f
cc_248 N_A_c_340_n N_B_c_529_n 2.15082e-19
cc_249 N_A_c_326_n N_B_c_502_n 0.00340226f
cc_250 N_A_c_332_n N_B_c_502_n 0.00192865f
cc_251 N_A_c_340_n N_B_c_502_n 6.44056e-19
cc_252 N_A_c_326_n N_B_c_514_n 5.44597e-19
cc_253 N_A_c_340_n N_Z_c_567_n 5.87699e-19
cc_254 N_A_XI28.X0_PGD N_Z_c_571_n 7.94638e-19
cc_255 N_A_c_332_n N_Z_c_571_n 0.00175701f
cc_256 N_A_c_340_n N_Z_c_571_n 0.00103031f
cc_257 N_BI_XI29.X0_CG N_AI_XI29.X0_PGD 9.47088e-19
cc_258 N_BI_c_418_n N_AI_XI29.X0_PGD 0.00133285f
cc_259 N_BI_c_399_n N_AI_c_463_n 8.39468e-19
cc_260 N_BI_c_392_n N_B_c_499_n 6.90199e-19
cc_261 N_BI_c_399_n N_B_c_501_n 0.00133142f
cc_262 N_BI_c_399_n N_B_c_537_n 5.44238e-19
cc_263 N_BI_c_428_p N_B_c_537_n 3.08318e-19
cc_264 N_BI_c_410_n N_B_c_512_n 0.00187472f
cc_265 N_BI_c_402_n N_B_c_512_n 0.00165773f
cc_266 N_BI_c_399_n N_B_c_541_n 4.56568e-19
cc_267 N_BI_c_418_n N_B_c_541_n 0.00266356f
cc_268 N_BI_c_419_n N_B_c_541_n 7.16621e-19
cc_269 N_BI_c_410_n N_B_c_529_n 4.62769e-19
cc_270 N_BI_c_418_n N_B_c_529_n 6.17967e-19
cc_271 N_BI_c_419_n N_B_c_529_n 0.00243633f
cc_272 N_BI_c_399_n N_B_c_502_n 0.00398399f
cc_273 N_BI_c_399_n N_B_c_548_n 3.07174e-19
cc_274 N_BI_c_402_n N_B_c_548_n 0.00126004f
cc_275 N_BI_c_440_p N_B_c_548_n 0.00342237f
cc_276 N_BI_c_399_n N_B_c_504_n 5.09978e-19
cc_277 N_BI_c_402_n N_B_c_504_n 9.4756e-19
cc_278 N_BI_c_428_p N_B_c_504_n 8.92139e-19
cc_279 N_BI_c_440_p N_B_c_554_n 0.00210118f
cc_280 N_BI_c_399_n N_B_c_505_n 0.00143025f
cc_281 N_BI_c_402_n N_B_c_505_n 9.46104e-19
cc_282 N_BI_c_399_n N_Z_c_571_n 0.00138952f
cc_283 N_BI_c_410_n N_Z_c_571_n 0.00141294f
cc_284 N_BI_c_418_n N_Z_c_571_n 8.66889e-19
cc_285 N_BI_c_419_n N_Z_c_571_n 8.66889e-19
cc_286 N_BI_c_402_n N_Z_c_571_n 0.00105522f
cc_287 N_BI_c_440_p N_Z_c_571_n 0.00212989f
cc_288 N_BI_c_428_p N_Z_c_571_n 0.00104995f
cc_289 N_AI_XI29.X0_PGD N_B_c_557_n 9.65637e-19
cc_290 N_AI_c_492_p N_B_c_537_n 2.15082e-19
cc_291 N_AI_XI29.X0_PGD N_B_c_541_n 0.00133285f
cc_292 N_AI_c_471_n N_B_c_541_n 2.15082e-19
cc_293 N_AI_c_492_p N_B_c_541_n 5.05931e-19
cc_294 N_AI_c_463_n N_B_c_502_n 4.67711e-19
cc_295 N_AI_XI29.X0_PGD N_Z_c_571_n 4.32017e-19
cc_296 N_B_c_537_n N_Z_c_571_n 0.00157325f
cc_297 N_B_c_512_n N_Z_c_571_n 0.00138952f
cc_298 N_B_c_529_n N_Z_c_571_n 8.66889e-19
cc_299 N_B_c_548_n N_Z_c_571_n 4.69528e-19
*
.ends
*
*
.subckt XOR3_HPNW12 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XOR3_N3
.ends
