* sclib_tigfet10_hpnw4_tt_0p70v_25c.sp
.subckt TIGFET_HPNW4 D PGD CG PGS S
xgate (D PGD CG PGS S) TIGFET nw=4
.ends
*
* File: G3_AND2_N1.pex.netlist
* Created: Wed Feb 23 10:37:48 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_AND2_N1_VSS 2 4 6 8 10 12 14 16 30 31 33 50 53 70 75 80 85 94 99
+ 108 109 113 114 119 125 127 132 133 134 136 Vss
c68 134 Vss 3.75522e-19
c69 133 Vss 3.62111e-19
c70 132 Vss 0.00361417f
c71 127 Vss 0.00255728f
c72 125 Vss 0.00548072f
c73 119 Vss 0.00398592f
c74 114 Vss 9.65205e-19
c75 113 Vss 0.00179171f
c76 109 Vss 8.2274e-19
c77 108 Vss 0.00426189f
c78 99 Vss 0.00393602f
c79 94 Vss 0.004332f
c80 85 Vss 7.10513e-22
c81 80 Vss 6.65776e-19
c82 75 Vss 3.89225e-19
c83 70 Vss 0.00133027f
c84 58 Vss 0.0299355f
c85 57 Vss 0.0299355f
c86 53 Vss 7.50699e-20
c87 51 Vss 0.0346861f
c88 50 Vss 0.0984533f
c89 42 Vss 0.105926f
c90 37 Vss 0.0688517f
c91 33 Vss 6.52493e-20
c92 31 Vss 0.0342473f
c93 30 Vss 0.064644f
c94 16 Vss 0.00266844f
c95 14 Vss 0.0828881f
c96 12 Vss 0.0825199f
c97 10 Vss 0.0830027f
c98 8 Vss 0.0831275f
c99 6 Vss 0.0832632f
c100 4 Vss 0.0828837f
c101 2 Vss 0.00266829f
r102 132 136 0.326018
r103 131 132 4.16786
r104 127 131 0.655813
r105 126 134 0.494161
r106 125 136 0.326018
r107 125 126 10.1279
r108 121 134 0.128424
r109 120 133 0.494161
r110 119 134 0.494161
r111 119 120 10.378
r112 115 133 0.128424
r113 113 133 0.494161
r114 113 114 4.37625
r115 108 114 0.668428
r116 107 109 0.6565
r117 107 108 10.093
r118 85 127 1.82344
r119 80 99 1.16709
r120 80 121 2.16729
r121 75 94 1.16709
r122 75 115 2.16729
r123 70 109 1.85991
r124 53 99 0.238214
r125 51 53 1.45875
r126 50 54 0.652036
r127 50 53 1.45875
r128 47 51 0.652036
r129 43 58 0.494161
r130 42 44 0.652036
r131 42 43 2.9175
r132 39 58 0.128424
r133 38 57 0.494161
r134 37 58 0.494161
r135 37 38 2.8008
r136 34 57 0.128424
r137 33 94 0.238214
r138 31 33 1.4004
r139 30 57 0.494161
r140 30 33 1.5171
r141 27 31 0.652036
r142 16 85 1.16709
r143 14 47 2.5674
r144 12 54 2.5674
r145 10 44 2.5674
r146 8 39 2.5674
r147 6 27 2.5674
r148 4 34 2.5674
r149 2 70 1.16709
.ends

.subckt PM_G3_AND2_N1_VDD 2 4 6 10 12 25 27 33 51 53 54 58 60 64 68 70 74 76 78
+ 79 85 94 Vss
c87 94 Vss 0.00555165f
c88 85 Vss 0.00507125f
c89 79 Vss 4.42156e-19
c90 76 Vss 5.947e-19
c91 74 Vss 0.00125165f
c92 70 Vss 0.00410186f
c93 68 Vss 0.0014864f
c94 64 Vss 0.0023623f
c95 60 Vss 0.00679469f
c96 58 Vss 0.0016182f
c97 55 Vss 0.00207011f
c98 54 Vss 0.0101277f
c99 53 Vss 0.0036687f
c100 51 Vss 0.00587536f
c101 33 Vss 0.0347789f
c102 32 Vss 0.101192f
c103 27 Vss 0.183894f
c104 25 Vss 0.0364084f
c105 12 Vss 0.0842982f
c106 10 Vss 0.0825186f
c107 6 Vss 0.00153036f
c108 4 Vss 0.00221866f
c109 2 Vss 0.0976708f
r110 74 94 1.16709
r111 72 74 2.16729
r112 71 79 0.494161
r113 70 72 0.652036
r114 70 71 7.46046
r115 66 79 0.128424
r116 66 68 4.83471
r117 64 85 1.16709
r118 62 64 3.66771
r119 61 78 0.386734
r120 60 79 0.494161
r121 60 61 13.0037
r122 56 76 0.18826
r123 56 58 1.82344
r124 54 62 0.652036
r125 54 55 10.0862
r126 53 78 0.284962
r127 52 76 0.427332
r128 52 53 3.07105
r129 51 76 0.427332
r130 50 55 0.671696
r131 50 51 7.86189
r132 35 94 0.238214
r133 33 35 1.45875
r134 32 36 0.652036
r135 32 35 1.45875
r136 29 33 0.652036
r137 27 85 0.50025
r138 25 27 5.11257
r139 22 25 0.652541
r140 12 36 2.5674
r141 10 29 2.5674
r142 6 68 1.16709
r143 4 58 1.16709
r144 2 22 3.2676
.ends

.subckt PM_G3_AND2_N1_A 2 4 10 13 18 21 26 31 Vss
c25 31 Vss 0.00351715f
c26 26 Vss 0.00299969f
c27 18 Vss 8.55683e-19
c28 13 Vss 0.0576606f
c29 2 Vss 0.0575116f
r30 23 31 1.16709
r31 21 23 2.12561
r32 18 26 1.16709
r33 18 21 2.70911
r34 13 31 0.50025
r35 10 26 0.50025
r36 4 13 1.80885
r37 2 10 1.80885
.ends

.subckt PM_G3_AND2_N1_NET1 2 4 8 10 21 24 27 45 53 66 70 Vss
c51 70 Vss 0.00676771f
c52 66 Vss 0.00607266f
c53 53 Vss 0.00254578f
c54 45 Vss 0.00159242f
c55 27 Vss 1.04894e-19
c56 24 Vss 0.225594f
c57 21 Vss 0.0713786f
c58 19 Vss 0.0247918f
c59 10 Vss 0.0847975f
c60 4 Vss 0.00148239f
c61 2 Vss 0.00144265f
r62 70 74 0.652036
r63 53 66 1.16709
r64 53 74 3.66771
r65 48 70 8.04396
r66 48 50 6.4185
r67 45 48 2.75079
r68 27 66 0.0476429
r69 25 27 0.326018
r70 25 27 0.1167
r71 24 28 0.652036
r72 24 27 6.7686
r73 21 66 0.357321
r74 19 27 0.326018
r75 19 21 0.40845
r76 10 28 2.5674
r77 8 21 2.15895
r78 4 50 1.16709
r79 2 45 1.16709
.ends

.subckt PM_G3_AND2_N1_B 2 4 10 11 14 18 21 Vss
c26 21 Vss 5.0923e-19
c27 14 Vss 0.148163f
c28 11 Vss 0.0348321f
c29 10 Vss 0.287297f
c30 2 Vss 0.172263f
r31 18 21 0.0364688
r32 14 21 1.16709
r33 12 14 2.8008
r34 10 12 0.652036
r35 10 11 8.92755
r36 7 11 0.652036
r37 4 14 3.0342
r38 2 7 5.835
.ends

.subckt PM_G3_AND2_N1_Z 2 16 19 Vss
c11 2 Vss 0.00148239f
r12 16 19 0.0364688
r13 2 19 1.16709
.ends

.subckt G3_AND2_N1  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI7.X0 N_NET1_XI7.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_B_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW4
XI8.X0 N_NET1_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI9.X0 N_NET1_XI8.X0_D N_VSS_XI9.X0_PGD N_B_XI9.X0_CG N_VSS_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW4
XI2.X0 N_Z_XI2.X0_D N_VSS_XI2.X0_PGD N_NET1_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW4
XI1.X0 N_Z_XI2.X0_D N_VDD_XI1.X0_PGD N_NET1_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
*
x_PM_G3_AND2_N1_VSS N_VSS_XI7.X0_S N_VSS_XI8.X0_PGD N_VSS_XI8.X0_PGS
+ N_VSS_XI9.X0_PGD N_VSS_XI9.X0_PGS N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI1.X0_S N_VSS_c_13_p N_VSS_c_14_p N_VSS_c_42_p N_VSS_c_2_p N_VSS_c_49_p
+ N_VSS_c_4_p N_VSS_c_7_p N_VSS_c_23_p N_VSS_c_65_p N_VSS_c_8_p N_VSS_c_25_p
+ N_VSS_c_5_p N_VSS_c_6_p N_VSS_c_17_p N_VSS_c_10_p N_VSS_c_18_p N_VSS_c_30_p
+ N_VSS_c_68_p N_VSS_c_33_p N_VSS_c_19_p N_VSS_c_31_p VSS Vss PM_G3_AND2_N1_VSS
x_PM_G3_AND2_N1_VDD N_VDD_XI7.X0_PGD N_VDD_XI8.X0_S N_VDD_XI9.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_c_143_p N_VDD_c_128_p N_VDD_c_70_n
+ N_VDD_c_71_n N_VDD_c_75_n N_VDD_c_79_n N_VDD_c_80_n N_VDD_c_81_n N_VDD_c_116_p
+ N_VDD_c_88_n N_VDD_c_94_n N_VDD_c_100_n N_VDD_c_102_n VDD N_VDD_c_103_n
+ N_VDD_c_113_p N_VDD_c_104_n Vss PM_G3_AND2_N1_VDD
x_PM_G3_AND2_N1_A N_A_XI7.X0_CG N_A_XI8.X0_CG N_A_c_164_n N_A_c_156_n
+ N_A_c_157_n A N_A_c_167_n N_A_c_160_n Vss PM_G3_AND2_N1_A
x_PM_G3_AND2_N1_NET1 N_NET1_XI7.X0_D N_NET1_XI8.X0_D N_NET1_XI2.X0_CG
+ N_NET1_XI1.X0_CG N_NET1_c_183_n N_NET1_c_184_n N_NET1_c_185_n N_NET1_c_187_n
+ N_NET1_c_190_n N_NET1_c_193_n N_NET1_c_195_n Vss PM_G3_AND2_N1_NET1
x_PM_G3_AND2_N1_B N_B_XI7.X0_PGS N_B_XI9.X0_CG N_B_c_232_n N_B_c_234_n
+ N_B_c_239_n B N_B_c_242_n Vss PM_G3_AND2_N1_B
x_PM_G3_AND2_N1_Z N_Z_XI2.X0_D Z N_Z_c_260_n Vss PM_G3_AND2_N1_Z
cc_1 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.0016786f
cc_2 N_VSS_c_2_p N_VDD_c_70_n 0.0016786f
cc_3 N_VSS_XI7.X0_S N_VDD_c_71_n 9.73142e-19
cc_4 N_VSS_c_4_p N_VDD_c_71_n 0.0016649f
cc_5 N_VSS_c_5_p N_VDD_c_71_n 0.00583639f
cc_6 N_VSS_c_6_p N_VDD_c_71_n 0.00213268f
cc_7 N_VSS_c_7_p N_VDD_c_75_n 9.61646e-19
cc_8 N_VSS_c_8_p N_VDD_c_75_n 4.3619e-19
cc_9 N_VSS_c_5_p N_VDD_c_75_n 0.00351219f
cc_10 N_VSS_c_10_p N_VDD_c_75_n 0.00128683f
cc_11 N_VSS_c_4_p N_VDD_c_79_n 0.00221042f
cc_12 N_VSS_c_4_p N_VDD_c_80_n 7.48389e-19
cc_13 N_VSS_c_13_p N_VDD_c_81_n 0.00144388f
cc_14 N_VSS_c_14_p N_VDD_c_81_n 2.81922e-19
cc_15 N_VSS_c_7_p N_VDD_c_81_n 0.00161703f
cc_16 N_VSS_c_8_p N_VDD_c_81_n 2.03837e-19
cc_17 N_VSS_c_17_p N_VDD_c_81_n 0.00338232f
cc_18 N_VSS_c_18_p N_VDD_c_81_n 0.00635521f
cc_19 N_VSS_c_19_p N_VDD_c_81_n 7.61747e-19
cc_20 N_VSS_XI9.X0_PGS N_VDD_c_88_n 2.28184e-19
cc_21 N_VSS_XI2.X0_PGS N_VDD_c_88_n 2.56778e-19
cc_22 N_VSS_c_7_p N_VDD_c_88_n 5.65664e-19
cc_23 N_VSS_c_23_p N_VDD_c_88_n 0.00181281f
cc_24 N_VSS_c_8_p N_VDD_c_88_n 2.30125e-19
cc_25 N_VSS_c_25_p N_VDD_c_88_n 9.55109e-19
cc_26 N_VSS_c_2_p N_VDD_c_94_n 4.8598e-19
cc_27 N_VSS_c_23_p N_VDD_c_94_n 0.00161703f
cc_28 N_VSS_c_25_p N_VDD_c_94_n 2.03837e-19
cc_29 N_VSS_c_18_p N_VDD_c_94_n 0.00145178f
cc_30 N_VSS_c_30_p N_VDD_c_94_n 0.00590089f
cc_31 N_VSS_c_31_p N_VDD_c_94_n 7.74609e-19
cc_32 N_VSS_c_23_p N_VDD_c_100_n 8.94411e-19
cc_33 N_VSS_c_33_p N_VDD_c_100_n 3.85245e-19
cc_34 N_VSS_c_5_p N_VDD_c_102_n 0.00104993f
cc_35 N_VSS_c_18_p N_VDD_c_103_n 0.00119068f
cc_36 N_VSS_c_23_p N_VDD_c_104_n 3.48267e-19
cc_37 N_VSS_c_25_p N_VDD_c_104_n 8.0279e-19
cc_38 N_VSS_c_8_p N_A_c_156_n 0.00234241f
cc_39 N_VSS_c_7_p N_A_c_157_n 8.12473e-19
cc_40 N_VSS_c_8_p N_A_c_157_n 5.42695e-19
cc_41 N_VSS_c_5_p N_A_c_157_n 6.55807e-19
cc_42 N_VSS_c_42_p N_A_c_160_n 7.84334e-19
cc_43 N_VSS_c_7_p N_A_c_160_n 4.56568e-19
cc_44 N_VSS_c_8_p N_A_c_160_n 0.00184767f
cc_45 N_VSS_XI7.X0_S N_NET1_XI7.X0_D 3.43419e-19
cc_46 N_VSS_c_4_p N_NET1_XI7.X0_D 3.48267e-19
cc_47 N_VSS_c_25_p N_NET1_c_183_n 0.00413078f
cc_48 N_VSS_XI2.X0_PGD N_NET1_c_184_n 4.20799e-19
cc_49 N_VSS_c_49_p N_NET1_c_185_n 9.28737e-19
cc_50 N_VSS_c_25_p N_NET1_c_185_n 2.03369e-19
cc_51 N_VSS_XI7.X0_S N_NET1_c_187_n 3.48267e-19
cc_52 N_VSS_c_4_p N_NET1_c_187_n 8.46599e-19
cc_53 N_VSS_c_5_p N_NET1_c_187_n 2.07501e-19
cc_54 N_VSS_c_23_p N_NET1_c_190_n 0.00125323f
cc_55 N_VSS_c_25_p N_NET1_c_190_n 4.64764e-19
cc_56 N_VSS_c_5_p N_NET1_c_190_n 3.39684e-19
cc_57 N_VSS_c_23_p N_NET1_c_193_n 4.56568e-19
cc_58 N_VSS_c_25_p N_NET1_c_193_n 6.1245e-19
cc_59 N_VSS_c_5_p N_NET1_c_195_n 2.06399e-19
cc_60 N_VSS_c_18_p N_NET1_c_195_n 0.00149275f
cc_61 N_VSS_XI8.X0_PGD N_B_c_232_n 6.72196e-19
cc_62 N_VSS_XI9.X0_PGD N_B_c_232_n 6.72196e-19
cc_63 N_VSS_XI8.X0_PGS N_B_c_234_n 7.85613e-19
cc_64 N_VSS_XI1.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_65 N_VSS_c_65_p N_Z_XI2.X0_D 3.48267e-19
cc_66 N_VSS_c_65_p N_Z_c_260_n 5.37696e-19
cc_67 N_VSS_c_30_p N_Z_c_260_n 2.64173e-19
cc_68 N_VSS_c_68_p N_Z_c_260_n 2.7826e-19
cc_69 N_VDD_XI7.X0_PGD N_A_XI7.X0_CG 4.88425e-19
cc_70 N_VDD_c_79_n N_A_c_164_n 3.72495e-19
cc_71 N_VDD_c_71_n N_A_c_157_n 0.00273528f
cc_72 N_VDD_c_79_n N_A_c_157_n 7.03725e-19
cc_73 N_VDD_XI7.X0_PGD N_A_c_167_n 2.88617e-19
cc_74 N_VDD_c_71_n N_A_c_167_n 3.68786e-19
cc_75 N_VDD_c_79_n N_A_c_167_n 4.3265e-19
cc_76 N_VDD_c_113_p N_A_c_167_n 7.96439e-19
cc_77 N_VDD_c_71_n N_A_c_160_n 5.09899e-19
cc_78 N_VDD_c_79_n N_NET1_XI7.X0_D 9.18655e-19
cc_79 N_VDD_c_116_p N_NET1_XI7.X0_D 8.835e-19
cc_80 N_VDD_c_113_p N_NET1_XI7.X0_D 0.00132057f
cc_81 N_VDD_XI8.X0_S N_NET1_XI8.X0_D 3.43419e-19
cc_82 N_VDD_XI9.X0_S N_NET1_XI8.X0_D 3.43419e-19
cc_83 N_VDD_c_80_n N_NET1_XI8.X0_D 3.74351e-19
cc_84 N_VDD_c_81_n N_NET1_XI8.X0_D 3.7884e-19
cc_85 N_VDD_c_88_n N_NET1_XI8.X0_D 3.48267e-19
cc_86 N_VDD_c_104_n N_NET1_XI1.X0_CG 8.03148e-19
cc_87 N_VDD_XI1.X0_PGD N_NET1_c_184_n 4.25379e-19
cc_88 N_VDD_XI7.X0_PGD N_NET1_c_187_n 2.94751e-19
cc_89 N_VDD_XI8.X0_S N_NET1_c_187_n 3.48267e-19
cc_90 N_VDD_XI9.X0_S N_NET1_c_187_n 3.48267e-19
cc_91 N_VDD_c_128_p N_NET1_c_187_n 5.10453e-19
cc_92 N_VDD_c_71_n N_NET1_c_187_n 6.49505e-19
cc_93 N_VDD_c_79_n N_NET1_c_187_n 0.00151981f
cc_94 N_VDD_c_80_n N_NET1_c_187_n 8.1398e-19
cc_95 N_VDD_c_81_n N_NET1_c_187_n 5.36364e-19
cc_96 N_VDD_c_116_p N_NET1_c_187_n 0.00366419f
cc_97 N_VDD_c_88_n N_NET1_c_187_n 7.99681e-19
cc_98 N_VDD_c_113_p N_NET1_c_187_n 8.835e-19
cc_99 N_VDD_c_79_n N_NET1_c_195_n 3.89533e-19
cc_100 N_VDD_c_81_n N_NET1_c_195_n 3.69547e-19
cc_101 N_VDD_c_116_p N_NET1_c_195_n 4.83374e-19
cc_102 N_VDD_c_88_n N_NET1_c_195_n 4.34102e-19
cc_103 N_VDD_XI7.X0_PGD N_B_XI7.X0_PGS 0.00320719f
cc_104 N_VDD_c_71_n N_B_XI7.X0_PGS 6.17633e-19
cc_105 N_VDD_c_79_n N_B_XI7.X0_PGS 2.2956e-19
cc_106 N_VDD_c_143_p N_B_c_232_n 0.00973324f
cc_107 N_VDD_c_81_n N_B_c_239_n 4.48125e-19
cc_108 N_VDD_c_116_p N_B_c_239_n 4.13122e-19
cc_109 N_VDD_c_113_p N_B_c_239_n 0.00150022f
cc_110 N_VDD_c_81_n N_B_c_242_n 2.66883e-19
cc_111 N_VDD_c_116_p N_B_c_242_n 3.55986e-19
cc_112 N_VDD_c_113_p N_B_c_242_n 3.81676e-19
cc_113 N_VDD_XI9.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_114 N_VDD_c_88_n N_Z_XI2.X0_D 3.48267e-19
cc_115 N_VDD_c_94_n N_Z_XI2.X0_D 3.7884e-19
cc_116 N_VDD_XI9.X0_S N_Z_c_260_n 3.48267e-19
cc_117 N_VDD_c_88_n N_Z_c_260_n 7.06424e-19
cc_118 N_VDD_c_94_n N_Z_c_260_n 5.12447e-19
cc_119 N_A_c_157_n N_NET1_c_187_n 0.00751692f
cc_120 N_A_c_167_n N_NET1_c_187_n 9.57699e-19
cc_121 N_A_c_160_n N_NET1_c_187_n 9.18163e-19
cc_122 N_A_XI7.X0_CG N_B_XI7.X0_PGS 4.5346e-19
cc_123 N_A_c_167_n N_B_XI7.X0_PGS 5.70584e-19
cc_124 N_A_c_157_n N_B_c_232_n 2.1473e-19
cc_125 N_A_c_167_n N_B_c_232_n 0.0014179f
cc_126 N_A_c_160_n N_B_c_232_n 0.00112482f
cc_127 N_A_c_160_n N_B_c_239_n 9.27569e-19
cc_128 N_NET1_c_187_n N_B_c_232_n 7.63501e-19
cc_129 N_NET1_c_187_n N_B_c_239_n 9.91045e-19
cc_130 N_NET1_c_190_n N_B_c_239_n 3.63713e-19
cc_131 N_NET1_c_193_n N_B_c_239_n 0.00197331f
cc_132 N_NET1_c_187_n N_B_c_242_n 0.00142922f
cc_133 N_NET1_c_190_n N_B_c_242_n 3.90886e-19
cc_134 N_NET1_c_193_n N_B_c_242_n 3.48267e-19
*
.ends
*
*
.subckt AND2_HPNW4 A B Y VDD VSS
xgate (VSS VDD A B Y) G3_AND2_N1
.ends
*
* File: G2_AOI21_N1.pex.netlist
* Created: Mon Apr 11 11:24:15 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_AOI21_N1_VSS 2 4 6 8 19 25 38 43 48 57 66 67 69 77 78 79 83 84 86
+ 88 89 Vss
c53 89 Vss 4.28045e-19
c54 86 Vss 0.00420179f
c55 84 Vss 0.00142701f
c56 83 Vss 8.42815e-19
c57 79 Vss 0.00125695f
c58 78 Vss 4.66086e-19
c59 77 Vss 0.00243143f
c60 69 Vss 0.00100335f
c61 68 Vss 0.00135524f
c62 67 Vss 0.00884313f
c63 66 Vss 0.00244299f
c64 57 Vss 0.00663377f
c65 48 Vss 1.70165e-19
c66 43 Vss 0.00203396f
c67 38 Vss 0.00129403f
c68 25 Vss 0.0827803f
c69 19 Vss 0.034042f
c70 18 Vss 0.0688517f
c71 8 Vss 0.0810091f
c72 6 Vss 0.00226958f
c73 4 Vss 0.0797379f
c74 2 Vss 0.00290534f
r75 85 89 0.551426
r76 85 86 13.3371
r77 84 89 0.551426
r78 83 88 0.326149
r79 83 84 4.12618
r80 79 89 0.0828784
r81 77 86 0.652036
r82 77 78 4.33457
r83 73 78 0.652036
r84 67 88 0.326149
r85 67 68 15.1308
r86 66 69 0.655813
r87 65 68 0.652298
r88 65 66 4.12618
r89 48 79 1.82344
r90 43 57 1.16709
r91 43 73 2.16729
r92 38 69 1.82344
r93 25 57 0.238214
r94 23 25 2.04225
r95 20 23 0.0685365
r96 18 23 0.5835
r97 18 19 2.8008
r98 15 19 0.652036
r99 8 20 2.5674
r100 6 48 1.16709
r101 4 15 2.5674
r102 2 38 1.16709
.ends

.subckt PM_G2_AOI21_N1_VDD 2 4 6 8 10 45 46 48 50 54 56 57 58 63 65 67 68 74 Vss
c60 74 Vss 0.00498639f
c61 68 Vss 3.56526e-19
c62 65 Vss 0.00188744f
c63 63 Vss 0.00658029f
c64 58 Vss 0.00166035f
c65 57 Vss 6.17427e-19
c66 56 Vss 0.0030725f
c67 54 Vss 0.0015334f
c68 50 Vss 0.0128179f
c69 48 Vss 0.00148319f
c70 46 Vss 0.00118366f
c71 45 Vss 0.00509044f
c72 33 Vss 0.0307391f
c73 26 Vss 0.10055f
c74 22 Vss 0.0348457f
c75 21 Vss 0.0712517f
c76 10 Vss 0.00241752f
c77 8 Vss 0.0830779f
c78 6 Vss 0.0830019f
c79 4 Vss 0.00285737f
c80 2 Vss 0.0825892f
r81 64 68 0.551426
r82 64 65 4.16786
r83 63 68 0.551426
r84 62 63 13.2955
r85 58 68 0.0828784
r86 58 60 1.82344
r87 56 62 0.652298
r88 56 57 4.22534
r89 54 74 1.16709
r90 52 57 0.652298
r91 52 54 2.12561
r92 51 67 0.326018
r93 50 65 0.652036
r94 50 51 15.6711
r95 46 48 1.82344
r96 45 67 0.326018
r97 44 46 0.655813
r98 44 45 4.16786
r99 29 74 0.238214
r100 27 33 0.494161
r101 27 29 1.45875
r102 26 30 0.652036
r103 26 29 1.45875
r104 23 33 0.128424
r105 21 33 0.494161
r106 21 22 2.8008
r107 18 22 0.652036
r108 10 60 1.16709
r109 8 30 2.5674
r110 6 23 2.5674
r111 4 48 1.16709
r112 2 18 2.5674
.ends

.subckt PM_G2_AOI21_N1_B 2 4 20 23 29 Vss
c19 29 Vss 0.00607059f
c20 23 Vss 9.01834e-19
c21 20 Vss 0.0916059f
c22 16 Vss 0.0586024f
c23 4 Vss 0.0980254f
c24 2 Vss 0.320472f
r25 26 29 1.16709
r26 23 26 0.0833571
r27 18 20 2.04225
r28 16 29 0.197068
r29 13 16 1.2837
r30 10 20 0.0685365
r31 8 18 0.0685365
r32 7 13 0.0685365
r33 4 10 3.0342
r34 2 8 8.6358
r35 2 7 2.5674
.ends

.subckt PM_G2_AOI21_N1_C 2 4 6 17 24 28 31 35 38 42 45 58 Vss
c45 58 Vss 0.00118496f
c46 45 Vss 0.00482667f
c47 38 Vss 0.00276154f
c48 31 Vss 0.00515878f
c49 28 Vss 0.0945059f
c50 24 Vss 0.0559062f
c51 17 Vss 1.54762e-19
c52 6 Vss 0.178585f
c53 4 Vss 0.147123f
c54 2 Vss 0.0809403f
r55 54 58 0.652036
r56 38 58 5.16814
r57 38 42 0.0416786
r58 31 45 1.16709
r59 31 54 8.58579
r60 31 35 0.0416786
r61 26 28 2.04225
r62 24 45 0.197068
r63 21 24 1.2837
r64 18 28 0.0685365
r65 17 38 1.16709
r66 13 26 0.0685365
r67 13 17 2.8008
r68 10 21 0.0685365
r69 6 18 5.835
r70 4 17 3.0342
r71 2 10 2.5674
.ends

.subckt PM_G2_AOI21_N1_Z 2 4 30 33 Vss
c30 30 Vss 0.00225284f
c31 4 Vss 0.00143442f
c32 2 Vss 0.00153036f
r33 33 35 3.83443
r34 30 33 5.33486
r35 4 35 1.16709
r36 2 30 1.16709
.ends

.subckt PM_G2_AOI21_N1_A 2 4 10 11 13 14 15 20 24 28 31 Vss
c37 31 Vss 4.87906e-19
c38 28 Vss 4.59888e-19
c39 24 Vss 1.50097e-19
c40 20 Vss 0.0822806f
c41 18 Vss 0.0247918f
c42 15 Vss 0.032139f
c43 14 Vss 0.0725371f
c44 13 Vss 0.0312529f
c45 11 Vss 0.0345237f
c46 10 Vss 0.122163f
c47 2 Vss 0.188674f
r48 28 31 1.16709
r49 24 31 0.262036
r50 20 31 0.238214
r51 18 24 0.326018
r52 18 20 0.64185
r53 15 24 2.50905
r54 14 24 0.326018
r55 14 24 0.1167
r56 13 15 0.652036
r57 12 13 1.22535
r58 10 12 0.652036
r59 10 11 3.09255
r60 7 11 0.652036
r61 4 20 2.4507
r62 2 7 6.1851
.ends

.subckt G2_AOI21_N1  VSS VDD B C Z A
*
* A	A
* Z	Z
* C	C
* B	B
* VDD	VDD
* VSS	VSS
XI1.X0 N_Z_XI1.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_B_XI1.X0_PGS N_VSS_XI1.X0_S
+ TIGFET_HPNW4
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_C_XI6.X0_PGS N_VDD_XI6.X0_S
+ TIGFET_HPNW4
XI5.X0 N_Z_XI1.X0_D N_VDD_XI5.X0_PGD N_C_XI5.X0_CG N_VDD_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW4
XI7.X0 N_Z_XI6.X0_D N_VSS_XI7.X0_PGD N_A_XI7.X0_CG N_C_XI7.X0_PGS N_VDD_XI7.X0_S
+ TIGFET_HPNW4
*
x_PM_G2_AOI21_N1_VSS N_VSS_XI1.X0_S N_VSS_XI6.X0_PGD N_VSS_XI5.X0_S
+ N_VSS_XI7.X0_PGD N_VSS_c_3_p N_VSS_c_46_p N_VSS_c_2_p N_VSS_c_4_p N_VSS_c_8_p
+ N_VSS_c_20_p N_VSS_c_23_p N_VSS_c_9_p N_VSS_c_1_p N_VSS_c_5_p N_VSS_c_6_p
+ N_VSS_c_13_p N_VSS_c_10_p N_VSS_c_16_p N_VSS_c_17_p VSS N_VSS_c_18_p Vss
+ PM_G2_AOI21_N1_VSS
x_PM_G2_AOI21_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI6.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI5.X0_PGS N_VDD_XI7.X0_S N_VDD_c_89_p N_VDD_c_54_n N_VDD_c_55_n
+ N_VDD_c_56_n N_VDD_c_77_p N_VDD_c_60_n N_VDD_c_64_n N_VDD_c_65_n N_VDD_c_67_n
+ N_VDD_c_72_n VDD N_VDD_c_75_n N_VDD_c_78_p Vss PM_G2_AOI21_N1_VDD
x_PM_G2_AOI21_N1_B N_B_XI1.X0_PGS N_B_XI6.X0_CG N_B_c_122_p B N_B_c_119_n Vss
+ PM_G2_AOI21_N1_B
x_PM_G2_AOI21_N1_C N_C_XI6.X0_PGS N_C_XI5.X0_CG N_C_XI7.X0_PGS N_C_c_143_n
+ N_C_c_146_n N_C_c_147_n N_C_c_134_n C N_C_c_136_n C N_C_c_137_n N_C_c_140_n
+ Vss PM_G2_AOI21_N1_C
x_PM_G2_AOI21_N1_Z N_Z_XI1.X0_D N_Z_XI6.X0_D N_Z_c_182_n Z Vss PM_G2_AOI21_N1_Z
x_PM_G2_AOI21_N1_A N_A_XI1.X0_CG N_A_XI7.X0_CG N_A_c_208_n N_A_c_225_n
+ N_A_c_226_n N_A_c_209_n N_A_c_227_n N_A_c_211_n N_A_c_212_n A N_A_c_216_n Vss
+ PM_G2_AOI21_N1_A
cc_1 N_VSS_c_1_p N_VDD_c_54_n 4.93612e-19
cc_2 N_VSS_c_2_p N_VDD_c_55_n 9.30121e-19
cc_3 N_VSS_c_3_p N_VDD_c_56_n 0.0011834f
cc_4 N_VSS_c_4_p N_VDD_c_56_n 0.00161703f
cc_5 N_VSS_c_5_p N_VDD_c_56_n 0.00445263f
cc_6 N_VSS_c_6_p N_VDD_c_56_n 0.00169823f
cc_7 N_VSS_XI5.X0_S N_VDD_c_60_n 3.83684e-19
cc_8 N_VSS_c_8_p N_VDD_c_60_n 4.79306e-19
cc_9 N_VSS_c_9_p N_VDD_c_60_n 0.0035571f
cc_10 N_VSS_c_10_p N_VDD_c_60_n 0.00109026f
cc_11 N_VSS_c_9_p N_VDD_c_64_n 0.00162315f
cc_12 N_VSS_c_8_p N_VDD_c_65_n 2.13058e-19
cc_13 N_VSS_c_13_p N_VDD_c_65_n 5.33968e-19
cc_14 N_VSS_XI5.X0_S N_VDD_c_67_n 9.5668e-19
cc_15 N_VSS_c_8_p N_VDD_c_67_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_67_n 0.00300233f
cc_17 N_VSS_c_17_p N_VDD_c_67_n 0.00605714f
cc_18 N_VSS_c_18_p N_VDD_c_67_n 8.91588e-19
cc_19 N_VSS_c_4_p N_VDD_c_72_n 4.42697e-19
cc_20 N_VSS_c_20_p N_VDD_c_72_n 3.70842e-19
cc_21 N_VSS_c_17_p N_VDD_c_72_n 0.00278561f
cc_22 N_VSS_c_17_p N_VDD_c_75_n 9.45256e-19
cc_23 N_VSS_c_23_p B 3.22996e-19
cc_24 N_VSS_c_9_p B 3.31649e-19
cc_25 N_VSS_XI6.X0_PGD N_C_XI6.X0_PGS 0.00161425f
cc_26 N_VSS_c_4_p N_C_c_134_n 5.88052e-19
cc_27 N_VSS_c_17_p N_C_c_134_n 0.00138265f
cc_28 N_VSS_c_17_p N_C_c_136_n 3.65158e-19
cc_29 N_VSS_XI6.X0_PGD N_C_c_137_n 3.23173e-19
cc_30 N_VSS_c_4_p N_C_c_137_n 3.44698e-19
cc_31 N_VSS_c_20_p N_C_c_137_n 3.34921e-19
cc_32 N_VSS_c_9_p N_C_c_140_n 0.00303126f
cc_33 N_VSS_c_17_p N_C_c_140_n 3.90377e-19
cc_34 N_VSS_XI1.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_35 N_VSS_XI5.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_XI1.X0_D 3.48267e-19
cc_37 N_VSS_c_8_p N_Z_XI1.X0_D 3.48267e-19
cc_38 N_VSS_XI1.X0_S N_Z_c_182_n 3.48267e-19
cc_39 N_VSS_XI5.X0_S N_Z_c_182_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_182_n 5.69026e-19
cc_41 N_VSS_c_8_p N_Z_c_182_n 5.69026e-19
cc_42 N_VSS_c_9_p N_Z_c_182_n 4.18012e-19
cc_43 N_VSS_c_17_p N_Z_c_182_n 5.20852e-19
cc_44 N_VSS_XI6.X0_PGD N_A_c_208_n 7.38139e-19
cc_45 N_VSS_XI7.X0_PGD N_A_c_209_n 0.00160007f
cc_46 N_VSS_c_46_p N_A_c_209_n 3.07681e-19
cc_47 N_VSS_c_20_p N_A_c_211_n 0.00255152f
cc_48 N_VSS_c_46_p N_A_c_212_n 8.89952e-19
cc_49 N_VSS_c_20_p N_A_c_212_n 2.75949e-19
cc_50 N_VSS_c_4_p A 5.37794e-19
cc_51 N_VSS_c_20_p A 4.56568e-19
cc_52 N_VSS_c_4_p N_A_c_216_n 4.56568e-19
cc_53 N_VSS_c_20_p N_A_c_216_n 6.1245e-19
cc_54 N_VDD_XI1.X0_PGD N_B_XI1.X0_PGS 0.0015605f
cc_55 N_VDD_c_77_p B 5.21626e-19
cc_56 N_VDD_c_78_p B 3.48267e-19
cc_57 N_VDD_XI1.X0_PGD N_B_c_119_n 3.73456e-19
cc_58 N_VDD_c_77_p N_B_c_119_n 4.2695e-19
cc_59 N_VDD_c_78_p N_B_c_119_n 5.71625e-19
cc_60 N_VDD_c_78_p N_C_XI5.X0_CG 0.00117555f
cc_61 N_VDD_c_77_p N_C_c_143_n 4.85469e-19
cc_62 N_VDD_c_67_n N_C_c_143_n 5.82627e-19
cc_63 N_VDD_c_78_p N_C_c_143_n 0.00182135f
cc_64 N_VDD_c_56_n N_C_c_146_n 3.54083e-19
cc_65 N_VDD_XI5.X0_PGS N_C_c_147_n 7.91098e-19
cc_66 N_VDD_c_67_n N_C_c_147_n 4.33233e-19
cc_67 N_VDD_c_89_p N_C_c_134_n 3.48763e-19
cc_68 N_VDD_c_55_n N_C_c_134_n 3.25844e-19
cc_69 N_VDD_c_56_n N_C_c_134_n 0.00156477f
cc_70 N_VDD_c_56_n N_C_c_136_n 7.40864e-19
cc_71 N_VDD_c_77_p N_C_c_136_n 5.82566e-19
cc_72 N_VDD_c_67_n N_C_c_136_n 4.90875e-19
cc_73 N_VDD_c_78_p N_C_c_136_n 4.56568e-19
cc_74 N_VDD_c_89_p N_C_c_137_n 4.55865e-19
cc_75 N_VDD_c_56_n N_C_c_137_n 2.55177e-19
cc_76 N_VDD_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_77 N_VDD_XI7.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_78 N_VDD_c_55_n N_Z_XI6.X0_D 3.72199e-19
cc_79 N_VDD_c_56_n N_Z_XI6.X0_D 3.7884e-19
cc_80 N_VDD_c_65_n N_Z_XI6.X0_D 3.72199e-19
cc_81 N_VDD_XI6.X0_S N_Z_c_182_n 3.48267e-19
cc_82 N_VDD_XI7.X0_S N_Z_c_182_n 3.48267e-19
cc_83 N_VDD_c_55_n N_Z_c_182_n 5.68773e-19
cc_84 N_VDD_c_56_n N_Z_c_182_n 6.9352e-19
cc_85 N_VDD_c_65_n N_Z_c_182_n 7.77875e-19
cc_86 N_VDD_c_67_n N_Z_c_182_n 9.95668e-19
cc_87 N_VDD_XI1.X0_PGD N_A_c_208_n 6.1925e-19
cc_88 N_VDD_XI5.X0_PGD N_A_c_209_n 3.67852e-19
cc_89 N_VDD_c_67_n A 3.35548e-19
cc_90 N_VDD_c_56_n N_A_c_216_n 2.29043e-19
cc_91 N_VDD_c_67_n N_A_c_216_n 3.66936e-19
cc_92 N_B_c_122_p N_C_XI6.X0_PGS 0.00189436f
cc_93 N_B_XI1.X0_PGS N_C_XI5.X0_CG 2.46172e-19
cc_94 N_B_c_122_p N_C_XI7.X0_PGS 4.95875e-19
cc_95 N_B_c_122_p N_C_c_146_n 3.12087e-19
cc_96 N_B_XI1.X0_PGS N_Z_c_182_n 2.61881e-19
cc_97 N_B_XI1.X0_PGS N_A_XI1.X0_CG 0.00900711f
cc_98 N_B_c_119_n N_A_XI1.X0_CG 0.00150571f
cc_99 N_B_c_122_p N_A_c_225_n 0.00163406f
cc_100 N_B_XI1.X0_PGS N_A_c_226_n 6.07734e-19
cc_101 N_B_c_122_p N_A_c_227_n 0.00136506f
cc_102 N_B_c_122_p N_A_c_216_n 2.87722e-19
cc_103 N_C_c_143_n N_Z_c_182_n 9.29334e-19
cc_104 N_C_c_134_n N_Z_c_182_n 0.00223036f
cc_105 N_C_c_136_n N_Z_c_182_n 0.00299789f
cc_106 N_C_c_140_n N_Z_c_182_n 2.70867e-19
cc_107 N_C_XI5.X0_CG N_A_XI1.X0_CG 5.49495e-19
cc_108 N_C_c_143_n N_A_XI1.X0_CG 5.65259e-19
cc_109 N_C_XI7.X0_PGS N_A_c_208_n 8.10159e-19
cc_110 N_C_c_147_n N_A_c_208_n 0.00121323f
cc_111 N_C_XI7.X0_PGS N_A_c_211_n 5.00154e-19
cc_112 N_C_c_143_n N_A_c_212_n 9.55393e-19
cc_113 N_C_c_143_n A 4.56568e-19
cc_114 N_C_c_136_n A 6.2998e-19
cc_115 N_C_XI7.X0_PGS N_A_c_216_n 0.00570455f
cc_116 N_C_c_143_n N_A_c_216_n 8.77002e-19
cc_117 N_C_c_147_n N_A_c_216_n 0.00119367f
cc_118 N_C_c_136_n N_A_c_216_n 4.56568e-19
cc_119 N_Z_c_182_n N_A_XI1.X0_CG 5.75111e-19
cc_120 N_Z_c_182_n N_A_c_208_n 4.34888e-19
cc_121 N_Z_c_182_n A 0.0015179f
cc_122 N_Z_c_182_n N_A_c_216_n 8.99071e-19
*
.ends
*
*
.subckt AOI21_HPNW4 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 B0 Y A0) G2_AOI21_N1
.ends
*
* File: G2_BUF1_N1.pex.netlist
* Created: Wed Mar  2 15:26:00 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_BUF1_N1_VDD 2 4 7 11 28 32 52 56 58 59 63 67 69 73 77 90 95 Vss
c58 95 Vss 0.00471589f
c59 90 Vss 0.0048335f
c60 80 Vss 7.0893e-19
c61 79 Vss 7.0893e-19
c62 77 Vss 0.00107913f
c63 73 Vss 0.00106523f
c64 70 Vss 0.00175834f
c65 69 Vss 0.00726612f
c66 67 Vss 0.00110053f
c67 63 Vss 0.00110053f
c68 60 Vss 0.00175834f
c69 59 Vss 0.00712138f
c70 58 Vss 0.00330526f
c71 56 Vss 0.00424287f
c72 52 Vss 0.00330526f
c73 32 Vss 0.0346129f
c74 31 Vss 0.101192f
c75 28 Vss 0.0346129f
c76 27 Vss 0.101192f
c77 11 Vss 0.16682f
c78 7 Vss 0.16682f
c79 4 Vss 0.00203161f
c80 2 Vss 0.00233151f
r81 77 95 1.16709
r82 75 77 2.16729
r83 73 90 1.16709
r84 71 73 2.16729
r85 69 75 0.652036
r86 69 70 10.1279
r87 65 80 0.0828784
r88 65 67 1.82344
r89 61 79 0.0828784
r90 61 63 1.82344
r91 59 71 0.652036
r92 59 60 10.1279
r93 58 70 0.652036
r94 57 80 0.551426
r95 57 58 4.16786
r96 54 80 0.551426
r97 54 56 3.45932
r98 53 79 0.551426
r99 53 56 1.45875
r100 52 79 0.551426
r101 51 60 0.652036
r102 51 52 4.16786
r103 34 95 0.238214
r104 32 34 1.45875
r105 31 38 0.652036
r106 31 34 1.45875
r107 30 90 0.238214
r108 28 30 1.45875
r109 27 35 0.652036
r110 27 30 1.45875
r111 24 32 0.652036
r112 21 28 0.652036
r113 11 38 2.5674
r114 11 24 2.5674
r115 7 35 2.5674
r116 7 21 2.5674
r117 4 67 1.16709
r118 2 63 1.16709
.ends

.subckt PM_G2_BUF1_N1_VSS 3 7 10 12 27 28 31 32 52 57 62 67 72 77 97 98 99 100
+ 101 105 110 114 116 Vss
c60 118 Vss 6.78504e-19
c61 117 Vss 6.78504e-19
c62 116 Vss 0.00235663f
c63 114 Vss 0.00287691f
c64 110 Vss 0.00235663f
c65 105 Vss 9.66804e-19
c66 101 Vss 8.0746e-19
c67 100 Vss 5.83649e-19
c68 99 Vss 0.00631424f
c69 98 Vss 5.83649e-19
c70 97 Vss 0.00625937f
c71 77 Vss 0.00398915f
c72 72 Vss 0.00399741f
c73 67 Vss 1.62164e-19
c74 62 Vss 3.56438e-22
c75 57 Vss 8.13664e-19
c76 52 Vss 7.92706e-19
c77 34 Vss 1.28632e-19
c78 32 Vss 0.0341976f
c79 31 Vss 0.0984533f
c80 28 Vss 0.0341976f
c81 27 Vss 0.0984533f
c82 12 Vss 0.00237948f
c83 10 Vss 0.00207958f
c84 7 Vss 0.16682f
c85 3 Vss 0.16682f
r86 115 118 0.551426
r87 115 116 4.16786
r88 112 118 0.551426
r89 112 114 2.12561
r90 111 117 0.551426
r91 111 114 2.79246
r92 110 117 0.551426
r93 109 110 4.16786
r94 105 118 0.0828784
r95 101 117 0.0828784
r96 99 116 0.652036
r97 99 100 10.1279
r98 97 109 0.652036
r99 97 98 10.1279
r100 93 100 0.652036
r101 89 98 0.652036
r102 67 105 1.82344
r103 62 101 1.82344
r104 57 77 1.16709
r105 57 93 2.16729
r106 52 72 1.16709
r107 52 89 2.16729
r108 34 77 0.238214
r109 32 34 1.45875
r110 31 38 0.652036
r111 31 34 1.45875
r112 30 72 0.238214
r113 28 30 1.45875
r114 27 35 0.652036
r115 27 30 1.45875
r116 24 32 0.652036
r117 21 28 0.652036
r118 12 67 1.16709
r119 10 62 1.16709
r120 7 38 2.5674
r121 7 24 2.5674
r122 3 35 2.5674
r123 3 21 2.5674
.ends

.subckt PM_G2_BUF1_N1_A 2 4 9 12 22 25 28 Vss
c18 28 Vss 0.00276471f
c19 25 Vss 3.55586e-19
c20 12 Vss 0.20721f
c21 9 Vss 0.0715834f
c22 7 Vss 0.0247918f
c23 4 Vss 0.0847975f
r24 25 28 1.16709
r25 22 25 0.0795682
r26 15 28 0.0476429
r27 13 15 0.326018
r28 13 15 0.1167
r29 12 16 0.652036
r30 12 15 6.7686
r31 9 28 0.357321
r32 7 15 0.326018
r33 7 9 0.40845
r34 4 16 2.5674
r35 2 9 2.15895
.ends

.subckt PM_G2_BUF1_N1_Z 2 19 Vss
c15 19 Vss 2.80869e-19
c16 2 Vss 0.00176567f
r17 16 19 0.0364688
r18 2 16 1.16709
.ends

.subckt PM_G2_BUF1_N1_NET17 2 4 6 18 36 41 50 58 Vss
c37 58 Vss 5.85801e-19
c38 50 Vss 0.00307045f
c39 41 Vss 0.0013766f
c40 36 Vss 0.00137137f
c41 22 Vss 0.0247918f
c42 19 Vss 0.0295882f
c43 18 Vss 0.176231f
c44 6 Vss 0.0715834f
c45 4 Vss 0.00176567f
c46 2 Vss 0.0847975f
r47 54 58 0.653045
r48 41 50 1.16709
r49 41 58 2.1395
r50 36 54 3.45932
r51 28 50 0.0476429
r52 26 50 0.357321
r53 22 28 0.326018
r54 22 26 0.40845
r55 19 28 6.7686
r56 18 28 0.326018
r57 18 28 0.1167
r58 15 19 0.652036
r59 6 26 2.15895
r60 4 36 1.16709
r61 2 15 2.5674
.ends

.subckt G2_BUF1_N1  VDD VSS A Z
*
* Z	Z
* A	A
* VSS	VSS
* VDD	VDD
XI3.X0 N_Z_XI3.X0_D N_VSS_XI3.X0_PGD N_NET17_XI3.X0_CG N_VSS_XI3.X0_PGD
+ N_VDD_XI3.X0_S TIGFET_HPNW4
XI2.X0 N_NET17_XI2.X0_D N_VSS_XI2.X0_PGD N_A_XI2.X0_CG N_VSS_XI2.X0_PGD
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI0.X0 N_Z_XI3.X0_D N_VDD_XI0.X0_PGD N_NET17_XI0.X0_CG N_VDD_XI0.X0_PGD
+ N_VSS_XI0.X0_S TIGFET_HPNW4
XI1.X0 N_NET17_XI2.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW4
*
x_PM_G2_BUF1_N1_VDD N_VDD_XI3.X0_S N_VDD_XI2.X0_S N_VDD_XI0.X0_PGD
+ N_VDD_XI1.X0_PGD N_VDD_c_3_p N_VDD_c_6_p N_VDD_c_9_p VDD N_VDD_c_13_p
+ N_VDD_c_4_p N_VDD_c_38_p N_VDD_c_43_p N_VDD_c_7_p N_VDD_c_11_p N_VDD_c_15_p
+ N_VDD_c_12_p N_VDD_c_16_p Vss PM_G2_BUF1_N1_VDD
x_PM_G2_BUF1_N1_VSS N_VSS_XI3.X0_PGD N_VSS_XI2.X0_PGD N_VSS_XI0.X0_S
+ N_VSS_XI1.X0_S N_VSS_c_61_n N_VSS_c_63_n N_VSS_c_64_n N_VSS_c_66_n
+ N_VSS_c_67_n N_VSS_c_71_n N_VSS_c_101_p N_VSS_c_110_p N_VSS_c_75_n
+ N_VSS_c_79_n N_VSS_c_83_n N_VSS_c_84_n N_VSS_c_85_n N_VSS_c_86_n N_VSS_c_104_p
+ N_VSS_c_112_p N_VSS_c_87_n VSS N_VSS_c_88_n Vss PM_G2_BUF1_N1_VSS
x_PM_G2_BUF1_N1_A N_A_XI2.X0_CG N_A_XI1.X0_CG N_A_c_124_n N_A_c_120_n A
+ N_A_c_122_n N_A_c_123_n Vss PM_G2_BUF1_N1_A
x_PM_G2_BUF1_N1_Z N_Z_XI3.X0_D Z Vss PM_G2_BUF1_N1_Z
x_PM_G2_BUF1_N1_NET17 N_NET17_XI3.X0_CG N_NET17_XI2.X0_D N_NET17_XI0.X0_CG
+ N_NET17_c_155_n N_NET17_c_157_n N_NET17_c_160_n N_NET17_c_164_n
+ N_NET17_c_168_n Vss PM_G2_BUF1_N1_NET17
cc_1 N_VDD_XI0.X0_PGD N_VSS_XI3.X0_PGD 0.00173038f
cc_2 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00173038f
cc_3 N_VDD_c_3_p N_VSS_c_61_n 0.00173038f
cc_4 N_VDD_c_4_p N_VSS_c_61_n 2.91357e-19
cc_5 N_VDD_c_4_p N_VSS_c_63_n 3.24852e-19
cc_6 N_VDD_c_6_p N_VSS_c_64_n 0.00173038f
cc_7 N_VDD_c_7_p N_VSS_c_64_n 2.91357e-19
cc_8 N_VDD_c_7_p N_VSS_c_66_n 3.24852e-19
cc_9 N_VDD_c_9_p N_VSS_c_67_n 8.69498e-19
cc_10 N_VDD_c_4_p N_VSS_c_67_n 0.00141228f
cc_11 N_VDD_c_11_p N_VSS_c_67_n 0.00106872f
cc_12 N_VDD_c_12_p N_VSS_c_67_n 3.48267e-19
cc_13 N_VDD_c_13_p N_VSS_c_71_n 8.69498e-19
cc_14 N_VDD_c_7_p N_VSS_c_71_n 0.00141228f
cc_15 N_VDD_c_15_p N_VSS_c_71_n 0.00106872f
cc_16 N_VDD_c_16_p N_VSS_c_71_n 3.48267e-19
cc_17 N_VDD_c_9_p N_VSS_c_75_n 3.66936e-19
cc_18 N_VDD_c_4_p N_VSS_c_75_n 0.00112249f
cc_19 N_VDD_c_11_p N_VSS_c_75_n 3.99794e-19
cc_20 N_VDD_c_12_p N_VSS_c_75_n 8.09245e-19
cc_21 N_VDD_c_13_p N_VSS_c_79_n 3.66936e-19
cc_22 N_VDD_c_7_p N_VSS_c_79_n 0.00112249f
cc_23 N_VDD_c_15_p N_VSS_c_79_n 3.99794e-19
cc_24 N_VDD_c_16_p N_VSS_c_79_n 8.09245e-19
cc_25 N_VDD_c_4_p N_VSS_c_83_n 0.00554293f
cc_26 N_VDD_c_4_p N_VSS_c_84_n 0.0017359f
cc_27 N_VDD_c_7_p N_VSS_c_85_n 0.00562924f
cc_28 N_VDD_c_7_p N_VSS_c_86_n 0.0017359f
cc_29 N_VDD_c_11_p N_VSS_c_87_n 3.85245e-19
cc_30 N_VDD_c_15_p N_VSS_c_88_n 3.85245e-19
cc_31 N_VDD_c_16_p N_A_XI1.X0_CG 0.00254294f
cc_32 N_VDD_XI0.X0_PGD N_A_c_120_n 4.08785e-19
cc_33 N_VDD_XI1.X0_PGD N_A_c_120_n 4.04053e-19
cc_34 VDD N_A_c_122_n 5.94555e-19
cc_35 VDD N_A_c_123_n 4.56718e-19
cc_36 N_VDD_XI3.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_37 N_VDD_c_4_p N_Z_XI3.X0_D 3.7884e-19
cc_38 N_VDD_c_38_p N_Z_XI3.X0_D 3.72199e-19
cc_39 N_VDD_XI3.X0_S Z 3.48267e-19
cc_40 N_VDD_c_4_p Z 5.12447e-19
cc_41 N_VDD_c_38_p Z 7.4527e-19
cc_42 N_VDD_XI2.X0_S N_NET17_XI2.X0_D 3.43419e-19
cc_43 N_VDD_c_43_p N_NET17_XI2.X0_D 3.72199e-19
cc_44 N_VDD_c_12_p N_NET17_XI0.X0_CG 0.0023817f
cc_45 N_VDD_XI0.X0_PGD N_NET17_c_155_n 4.04053e-19
cc_46 N_VDD_XI1.X0_PGD N_NET17_c_155_n 4.08785e-19
cc_47 N_VDD_XI2.X0_S N_NET17_c_157_n 3.48267e-19
cc_48 N_VDD_c_43_p N_NET17_c_157_n 8.0086e-19
cc_49 N_VDD_c_7_p N_NET17_c_157_n 5.01863e-19
cc_50 N_VDD_c_11_p N_NET17_c_160_n 6.85072e-19
cc_51 N_VDD_c_15_p N_NET17_c_160_n 3.98507e-19
cc_52 N_VDD_c_12_p N_NET17_c_160_n 4.99367e-19
cc_53 N_VDD_c_16_p N_NET17_c_160_n 3.0441e-19
cc_54 N_VDD_c_11_p N_NET17_c_164_n 4.85469e-19
cc_55 N_VDD_c_15_p N_NET17_c_164_n 3.00204e-19
cc_56 N_VDD_c_12_p N_NET17_c_164_n 0.0014909f
cc_57 N_VDD_c_16_p N_NET17_c_164_n 6.61247e-19
cc_58 VDD N_NET17_c_168_n 3.1911e-19
cc_59 N_VSS_c_79_n N_A_c_124_n 0.0023454f
cc_60 N_VSS_XI3.X0_PGD N_A_c_120_n 4.07282e-19
cc_61 N_VSS_XI2.X0_PGD N_A_c_120_n 3.99472e-19
cc_62 N_VSS_c_67_n N_A_c_122_n 2.85158e-19
cc_63 N_VSS_c_71_n N_A_c_122_n 5.53028e-19
cc_64 N_VSS_c_75_n N_A_c_122_n 3.0441e-19
cc_65 N_VSS_c_79_n N_A_c_122_n 4.99367e-19
cc_66 N_VSS_c_67_n N_A_c_123_n 2.82333e-19
cc_67 N_VSS_c_71_n N_A_c_123_n 4.56568e-19
cc_68 N_VSS_c_75_n N_A_c_123_n 6.61247e-19
cc_69 N_VSS_c_79_n N_A_c_123_n 0.0014909f
cc_70 N_VSS_XI0.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_71 N_VSS_c_101_p N_Z_XI3.X0_D 3.48267e-19
cc_72 N_VSS_XI0.X0_S Z 3.48267e-19
cc_73 N_VSS_c_101_p Z 4.99861e-19
cc_74 N_VSS_c_104_p Z 2.7826e-19
cc_75 N_VSS_c_75_n N_NET17_XI3.X0_CG 0.00250664f
cc_76 N_VSS_XI1.X0_S N_NET17_XI2.X0_D 3.43419e-19
cc_77 N_VSS_XI3.X0_PGD N_NET17_c_155_n 3.99472e-19
cc_78 N_VSS_XI2.X0_PGD N_NET17_c_155_n 4.07282e-19
cc_79 N_VSS_XI1.X0_S N_NET17_c_157_n 3.48267e-19
cc_80 N_VSS_c_110_p N_NET17_c_157_n 4.8288e-19
cc_81 N_VSS_c_85_n N_NET17_c_157_n 5.36354e-19
cc_82 N_VSS_c_112_p N_NET17_c_157_n 5.49885e-19
cc_83 VSS N_NET17_c_157_n 6.44069e-19
cc_84 N_VSS_c_83_n N_NET17_c_160_n 3.16821e-19
cc_85 N_VSS_c_85_n N_NET17_c_160_n 2.03753e-19
cc_86 VSS N_NET17_c_160_n 8.09756e-19
cc_87 N_VSS_c_83_n N_NET17_c_168_n 0.00101305f
cc_88 N_VSS_c_85_n N_NET17_c_168_n 5.70583e-19
cc_89 N_A_c_120_n N_NET17_c_155_n 0.00954069f
cc_90 N_A_c_122_n N_NET17_c_157_n 8.44937e-19
cc_91 N_Z_XI3.X0_D N_NET17_XI2.X0_D 2.56268e-19
cc_92 Z N_NET17_XI2.X0_D 3.17139e-19
cc_93 N_Z_XI3.X0_D N_NET17_c_157_n 3.17139e-19
cc_94 Z N_NET17_c_157_n 3.16516e-19
*
.ends
*
*
.subckt BUF1_HPNW4 A Y VDD VSS
xgate (VDD VSS A Y) G2_BUF1_N1
.ends
*
* File: G3_DFFQ1_N1.pex.netlist
* Created: Tue Apr  5 22:58:19 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_DFFQ1_N1_VSS 2 4 6 8 10 12 14 29 42 44 49 67 72 78 83 88 93 102
+ 111 116 125 126 127 128 132 137 142 148 154 156 161 163 165 166 167 Vss
c117 167 Vss 4.28045e-19
c118 166 Vss 3.75522e-19
c119 165 Vss 3.75522e-19
c120 164 Vss 6.13404e-19
c121 163 Vss 0.00437039f
c122 161 Vss 0.00140798f
c123 156 Vss 0.00134457f
c124 154 Vss 0.0025067f
c125 148 Vss 0.00439094f
c126 142 Vss 0.00297776f
c127 132 Vss 0.00193747f
c128 128 Vss 7.01403e-19
c129 127 Vss 8.12244e-19
c130 126 Vss 0.00567951f
c131 125 Vss 0.00148961f
c132 116 Vss 0.00596988f
c133 111 Vss 0.00418189f
c134 102 Vss 0.00407665f
c135 93 Vss 1.70165e-19
c136 88 Vss 0.00119073f
c137 83 Vss 5.15444e-19
c138 78 Vss 0.00173585f
c139 72 Vss 0.00866259f
c140 67 Vss 0.00134806f
c141 49 Vss 0.0560391f
c142 44 Vss 0.0560391f
c143 42 Vss 7.82991e-20
c144 29 Vss 0.0355813f
c145 28 Vss 0.101268f
c146 14 Vss 0.0832368f
c147 12 Vss 0.00370216f
c148 10 Vss 0.0027334f
c149 8 Vss 0.0822683f
c150 6 Vss 0.0792534f
c151 4 Vss 0.0793599f
c152 2 Vss 0.00198471f
r153 162 167 0.551426
r154 162 163 13.3371
r155 161 167 0.551426
r156 160 161 4.16786
r157 156 167 0.0828784
r158 155 166 0.494161
r159 154 163 0.652036
r160 154 155 4.37625
r161 150 166 0.128424
r162 149 165 0.494161
r163 148 160 0.652036
r164 148 149 10.1279
r165 144 165 0.128424
r166 143 164 0.494161
r167 142 166 0.494161
r168 142 143 7.46046
r169 138 164 0.128424
r170 132 164 0.494161
r171 132 137 1.00029
r172 126 165 0.494161
r173 126 127 15.8795
r174 125 128 0.655813
r175 124 127 0.652036
r176 124 125 4.16786
r177 93 156 1.82344
r178 88 116 1.16709
r179 88 150 2.16729
r180 83 111 1.16709
r181 83 144 2.16729
r182 78 138 4.83471
r183 75 137 1.29204
r184 72 102 1.16709
r185 72 75 12.4202
r186 67 128 1.82344
r187 49 116 0.197068
r188 46 49 1.2837
r189 42 111 0.197068
r190 42 44 1.2837
r191 38 46 0.0685365
r192 35 44 0.0685365
r193 31 102 0.0476429
r194 29 31 1.45875
r195 28 32 0.652036
r196 28 31 1.45875
r197 25 29 0.652036
r198 14 38 2.5674
r199 12 93 1.16709
r200 10 78 1.16709
r201 8 35 2.5674
r202 6 32 2.5674
r203 4 25 2.5674
r204 2 67 1.16709
.ends

.subckt PM_G3_DFFQ1_N1_CK 2 4 6 8 18 25 37 40 Vss
c31 40 Vss 0.00572916f
c32 37 Vss 3.65059e-19
c33 33 Vss 0.0299355f
c34 25 Vss 0.165118f
c35 18 Vss 0.186407f
c36 15 Vss 0.077884f
c37 13 Vss 0.0247918f
c38 6 Vss 0.441644f
c39 4 Vss 0.0840059f
r40 37 40 1.16709
r41 26 33 0.494161
r42 25 27 0.652036
r43 25 26 4.84305
r44 22 33 0.128424
r45 21 40 0.238214
r46 19 21 0.326018
r47 19 21 0.1167
r48 18 33 0.494161
r49 18 21 6.7686
r50 15 21 0.262036
r51 13 21 0.326018
r52 13 15 0.05835
r53 6 8 12.837
r54 6 27 2.5674
r55 4 22 2.5674
r56 2 15 2.50905
.ends

.subckt PM_G3_DFFQ1_N1_VDD 2 4 6 10 12 14 28 42 44 49 63 64 65 70 72 76 78 79 82
+ 84 86 91 93 95 96 98 99 100 102 104 113 118 Vss
c117 118 Vss 0.00660773f
c118 113 Vss 0.00546672f
c119 104 Vss 0.00477384f
c120 100 Vss 3.56526e-19
c121 99 Vss 2.39889e-19
c122 98 Vss 4.42156e-19
c123 96 Vss 0.00351049f
c124 95 Vss 5.22595e-19
c125 93 Vss 0.00279817f
c126 91 Vss 0.00684574f
c127 86 Vss 0.00166444f
c128 84 Vss 0.00296655f
c129 82 Vss 0.00146489f
c130 79 Vss 4.90412e-19
c131 78 Vss 0.00554983f
c132 76 Vss 5.91088e-19
c133 72 Vss 0.00336584f
c134 70 Vss 0.00240239f
c135 67 Vss 0.00178747f
c136 65 Vss 8.63831e-19
c137 64 Vss 0.00713032f
c138 63 Vss 0.00360153f
c139 49 Vss 0.0578141f
c140 44 Vss 0.0572437f
c141 42 Vss 7.44761e-20
c142 29 Vss 0.0373466f
c143 28 Vss 0.100964f
c144 14 Vss 0.00374907f
c145 12 Vss 0.0826302f
c146 10 Vss 0.0827668f
c147 6 Vss 0.00176834f
c148 4 Vss 0.0823731f
c149 2 Vss 0.0811326f
r150 95 104 1.16709
r151 95 96 0.470345
r152 93 102 0.326018
r153 92 100 0.551426
r154 92 93 4.16786
r155 91 100 0.551426
r156 90 91 13.3371
r157 86 100 0.0828784
r158 86 88 1.82344
r159 85 99 0.494161
r160 84 90 0.652036
r161 84 85 4.37625
r162 82 118 1.16709
r163 80 99 0.128424
r164 80 82 2.16729
r165 78 102 0.326018
r166 78 79 10.1279
r167 76 113 1.16709
r168 74 79 0.652036
r169 74 76 2.16729
r170 73 98 0.494161
r171 72 99 0.494161
r172 72 73 7.46046
r173 68 98 0.128424
r174 68 70 4.83471
r175 67 96 3.82922
r176 64 98 0.494161
r177 64 65 13.0037
r178 63 67 0.655813
r179 62 65 0.652036
r180 62 63 7.002
r181 49 118 0.197068
r182 46 49 1.2837
r183 42 113 0.197068
r184 42 44 1.2837
r185 38 46 0.0685365
r186 35 44 0.0685365
r187 31 104 0.0476429
r188 29 31 1.45875
r189 28 32 0.652036
r190 28 31 1.45875
r191 25 29 0.652036
r192 14 88 1.16709
r193 12 38 2.5674
r194 10 35 2.5674
r195 6 70 1.16709
r196 4 25 2.5674
r197 2 32 2.5674
.ends

.subckt PM_G3_DFFQ1_N1_CKN 2 6 8 18 28 33 50 Vss
c38 51 Vss 0.00127799f
c39 50 Vss 0.0053557f
c40 33 Vss 6.7412e-19
c41 28 Vss 0.00188103f
c42 18 Vss 8.89292e-19
c43 6 Vss 0.365937f
c44 2 Vss 0.00148239f
r45 50 51 14.6709
r46 46 51 0.652036
r47 33 50 0.531835
r48 28 46 4.00114
r49 18 33 1.16709
r50 8 18 6.4185
r51 6 18 6.4185
r52 2 28 1.16709
.ends

.subckt PM_G3_DFFQ1_N1_D 2 4 11 12 22 25 28 Vss
c27 28 Vss 0.00185315f
c28 25 Vss 4.49891e-19
c29 12 Vss 0.210787f
c30 11 Vss 2.35358e-19
c31 7 Vss 0.0247918f
c32 4 Vss 0.0830137f
c33 2 Vss 0.0713067f
r34 25 28 1.16709
r35 22 25 0.0364688
r36 15 28 0.0476429
r37 13 15 0.326018
r38 13 15 0.1167
r39 12 16 0.652036
r40 12 15 6.7686
r41 11 28 0.357321
r42 7 15 0.326018
r43 7 11 0.40845
r44 4 16 2.5674
r45 2 11 2.15895
.ends

.subckt PM_G3_DFFQ1_N1_X 2 4 8 17 20 23 35 39 41 47 Vss
c50 47 Vss 0.00138877f
c51 41 Vss 6.77172e-19
c52 39 Vss 0.0010541f
c53 35 Vss 0.00217231f
c54 23 Vss 7.53039e-20
c55 20 Vss 0.21062f
c56 17 Vss 0.0712602f
c57 15 Vss 0.0247918f
c58 8 Vss 0.0829593f
c59 2 Vss 0.00172036f
r60 44 47 1.16709
r61 41 44 2.08393
r62 37 39 4.33457
r63 36 41 0.0685365
r64 35 37 0.652036
r65 35 36 1.70882
r66 23 47 0.0476429
r67 21 23 0.326018
r68 21 23 0.1167
r69 20 24 0.652036
r70 20 23 6.7686
r71 17 47 0.357321
r72 15 23 0.326018
r73 15 17 0.40845
r74 8 24 2.5674
r75 4 17 2.15895
r76 2 39 1.16709
.ends

.subckt PM_G3_DFFQ1_N1_Q 2 16 Vss
c12 16 Vss 4.30842e-19
c13 2 Vss 0.00150258f
r14 16 19 0.0416786
r15 2 19 1.16709
.ends

.subckt G3_DFFQ1_N1  VSS CK VDD D Q
*
* Q	Q
* D	D
* VDD	VDD
* CK	CK
* VSS	VSS
XI1.X0 N_CKN_XI1.X0_D N_VDD_XI1.X0_PGD N_CK_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI2.X0 N_CKN_XI1.X0_D N_VSS_XI2.X0_PGD N_CK_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI5.X0 N_X_XI5.X0_D N_VSS_XI5.X0_PGD N_D_XI5.X0_CG N_CK_XI5.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI3.X0 N_Q_XI3.X0_D N_VDD_XI3.X0_PGD N_X_XI3.X0_CG N_CK_XI3.X0_PGS
+ N_VSS_XI3.X0_S TIGFET_HPNW4
XI4.X0 N_X_XI5.X0_D N_VDD_XI4.X0_PGD N_D_XI4.X0_CG N_CKN_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW4
XI0.X0 N_Q_XI3.X0_D N_VSS_XI0.X0_PGD N_X_XI0.X0_CG N_CKN_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW4
*
x_PM_G3_DFFQ1_N1_VSS N_VSS_XI1.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI5.X0_PGD N_VSS_XI3.X0_S N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_11_p
+ N_VSS_c_89_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_15_p N_VSS_c_3_p N_VSS_c_32_p
+ N_VSS_c_23_p N_VSS_c_33_p N_VSS_c_45_p N_VSS_c_20_p N_VSS_c_4_p N_VSS_c_34_p
+ N_VSS_c_16_p N_VSS_c_7_p N_VSS_c_22_p N_VSS_c_17_p N_VSS_c_85_p VSS
+ N_VSS_c_38_p N_VSS_c_29_p N_VSS_c_39_p N_VSS_c_48_p N_VSS_c_51_p N_VSS_c_52_p
+ N_VSS_c_30_p N_VSS_c_40_p N_VSS_c_53_p Vss PM_G3_DFFQ1_N1_VSS
x_PM_G3_DFFQ1_N1_CK N_CK_XI1.X0_CG N_CK_XI2.X0_CG N_CK_XI5.X0_PGS
+ N_CK_XI3.X0_PGS N_CK_c_122_n N_CK_c_123_n CK N_CK_c_129_p Vss
+ PM_G3_DFFQ1_N1_CK
x_PM_G3_DFFQ1_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI2.X0_S
+ N_VDD_XI3.X0_PGD N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_152_n N_VDD_c_250_p
+ N_VDD_c_153_n N_VDD_c_154_n N_VDD_c_155_n N_VDD_c_159_n N_VDD_c_163_n
+ N_VDD_c_164_n N_VDD_c_166_n N_VDD_c_172_n N_VDD_c_176_n N_VDD_c_182_n
+ N_VDD_c_183_n N_VDD_c_185_n N_VDD_c_188_n N_VDD_c_190_n N_VDD_c_195_n
+ N_VDD_c_199_n N_VDD_c_201_n N_VDD_c_203_n N_VDD_c_204_n N_VDD_c_205_n VDD
+ N_VDD_c_206_n N_VDD_c_208_n N_VDD_c_211_n Vss PM_G3_DFFQ1_N1_VDD
x_PM_G3_DFFQ1_N1_CKN N_CKN_XI1.X0_D N_CKN_XI4.X0_PGS N_CKN_XI0.X0_PGS
+ N_CKN_c_283_n N_CKN_c_268_n N_CKN_c_272_n N_CKN_c_274_n Vss PM_G3_DFFQ1_N1_CKN
x_PM_G3_DFFQ1_N1_D N_D_XI5.X0_CG N_D_XI4.X0_CG N_D_c_305_n N_D_c_306_n D
+ N_D_c_308_n N_D_c_312_n Vss PM_G3_DFFQ1_N1_D
x_PM_G3_DFFQ1_N1_X N_X_XI5.X0_D N_X_XI3.X0_CG N_X_XI0.X0_CG N_X_c_346_n
+ N_X_c_334_n N_X_c_354_n N_X_c_336_n N_X_c_337_n N_X_c_341_n N_X_c_343_n Vss
+ PM_G3_DFFQ1_N1_X
x_PM_G3_DFFQ1_N1_Q N_Q_XI3.X0_D Q Vss PM_G3_DFFQ1_N1_Q
cc_1 N_VSS_XI2.X0_PGS N_CK_XI5.X0_PGS 0.0029499f
cc_2 N_VSS_XI5.X0_PGD N_CK_XI5.X0_PGS 0.00158255f
cc_3 N_VSS_c_3_p N_CK_XI5.X0_PGS 8.20198e-19
cc_4 N_VSS_c_4_p N_CK_XI5.X0_PGS 4.62582e-19
cc_5 N_VSS_XI2.X0_PGD N_CK_c_122_n 4.16623e-19
cc_6 N_VSS_XI2.X0_PGS N_CK_c_123_n 4.26524e-19
cc_7 N_VSS_c_7_p CK 5.33707e-19
cc_8 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.00168612f
cc_9 N_VSS_XI0.X0_PGD N_VDD_XI3.X0_PGD 0.00189944f
cc_10 N_VSS_XI5.X0_PGD N_VDD_XI4.X0_PGD 0.00180681f
cc_11 N_VSS_c_11_p N_VDD_c_152_n 0.00168612f
cc_12 N_VSS_c_12_p N_VDD_c_153_n 0.00189944f
cc_13 N_VSS_c_13_p N_VDD_c_154_n 0.00180681f
cc_14 N_VSS_XI1.X0_S N_VDD_c_155_n 9.5668e-19
cc_15 N_VSS_c_15_p N_VDD_c_155_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_155_n 0.00321182f
cc_17 N_VSS_c_17_p N_VDD_c_155_n 0.00182807f
cc_18 N_VSS_c_15_p N_VDD_c_159_n 5.16845e-19
cc_19 N_VSS_c_3_p N_VDD_c_159_n 2.61925e-19
cc_20 N_VSS_c_20_p N_VDD_c_159_n 4.48125e-19
cc_21 N_VSS_c_7_p N_VDD_c_159_n 0.00922264f
cc_22 N_VSS_c_22_p N_VDD_c_163_n 0.00105444f
cc_23 N_VSS_c_23_p N_VDD_c_164_n 0.00239254f
cc_24 N_VSS_c_4_p N_VDD_c_164_n 9.55109e-19
cc_25 N_VSS_c_13_p N_VDD_c_166_n 2.43144e-19
cc_26 N_VSS_c_23_p N_VDD_c_166_n 0.00161703f
cc_27 N_VSS_c_4_p N_VDD_c_166_n 2.03837e-19
cc_28 N_VSS_c_7_p N_VDD_c_166_n 0.00131925f
cc_29 N_VSS_c_29_p N_VDD_c_166_n 0.00399563f
cc_30 N_VSS_c_30_p N_VDD_c_166_n 7.74609e-19
cc_31 N_VSS_c_3_p N_VDD_c_172_n 0.00179177f
cc_32 N_VSS_c_32_p N_VDD_c_172_n 3.92901e-19
cc_33 N_VSS_c_33_p N_VDD_c_172_n 8.51944e-19
cc_34 N_VSS_c_34_p N_VDD_c_172_n 3.99794e-19
cc_35 N_VSS_c_12_p N_VDD_c_176_n 3.37151e-19
cc_36 N_VSS_c_33_p N_VDD_c_176_n 0.00141228f
cc_37 N_VSS_c_34_p N_VDD_c_176_n 0.00112249f
cc_38 N_VSS_c_38_p N_VDD_c_176_n 0.00402042f
cc_39 N_VSS_c_39_p N_VDD_c_176_n 0.00326829f
cc_40 N_VSS_c_40_p N_VDD_c_176_n 7.74609e-19
cc_41 N_VSS_c_38_p N_VDD_c_182_n 0.00142104f
cc_42 N_VSS_c_23_p N_VDD_c_183_n 9.29543e-19
cc_43 N_VSS_c_4_p N_VDD_c_183_n 3.82294e-19
cc_44 N_VSS_XI4.X0_S N_VDD_c_185_n 3.7884e-19
cc_45 N_VSS_c_45_p N_VDD_c_185_n 4.73473e-19
cc_46 N_VSS_c_29_p N_VDD_c_185_n 0.00432522f
cc_47 N_VSS_c_45_p N_VDD_c_188_n 2.14355e-19
cc_48 N_VSS_c_48_p N_VDD_c_188_n 5.52785e-19
cc_49 N_VSS_XI4.X0_S N_VDD_c_190_n 9.5668e-19
cc_50 N_VSS_c_45_p N_VDD_c_190_n 0.00165395f
cc_51 N_VSS_c_51_p N_VDD_c_190_n 0.00302432f
cc_52 N_VSS_c_52_p N_VDD_c_190_n 0.00617602f
cc_53 N_VSS_c_53_p N_VDD_c_190_n 8.91588e-19
cc_54 N_VSS_c_33_p N_VDD_c_195_n 4.43871e-19
cc_55 N_VSS_c_34_p N_VDD_c_195_n 3.66936e-19
cc_56 N_VSS_c_39_p N_VDD_c_195_n 0.00106633f
cc_57 N_VSS_c_52_p N_VDD_c_195_n 0.00303537f
cc_58 N_VSS_c_3_p N_VDD_c_199_n 6.19689e-19
cc_59 N_VSS_c_20_p N_VDD_c_199_n 3.8721e-19
cc_60 N_VSS_c_15_p N_VDD_c_201_n 0.00303908f
cc_61 N_VSS_c_7_p N_VDD_c_201_n 2.94014e-19
cc_62 N_VSS_c_7_p N_VDD_c_203_n 0.00116322f
cc_63 N_VSS_c_29_p N_VDD_c_204_n 0.00102846f
cc_64 N_VSS_c_52_p N_VDD_c_205_n 0.00116512f
cc_65 N_VSS_c_3_p N_VDD_c_206_n 3.86162e-19
cc_66 N_VSS_c_20_p N_VDD_c_206_n 6.0892e-19
cc_67 N_VSS_c_3_p N_VDD_c_208_n 5.29489e-19
cc_68 N_VSS_c_33_p N_VDD_c_208_n 3.48267e-19
cc_69 N_VSS_c_34_p N_VDD_c_208_n 8.07896e-19
cc_70 N_VSS_c_23_p N_VDD_c_211_n 3.48267e-19
cc_71 N_VSS_c_4_p N_VDD_c_211_n 8.0279e-19
cc_72 N_VSS_XI1.X0_S N_CKN_XI1.X0_D 3.43419e-19
cc_73 N_VSS_c_15_p N_CKN_XI1.X0_D 3.48267e-19
cc_74 N_VSS_XI1.X0_S N_CKN_c_268_n 3.48267e-19
cc_75 N_VSS_c_15_p N_CKN_c_268_n 0.00105962f
cc_76 N_VSS_c_3_p N_CKN_c_268_n 7.53164e-19
cc_77 N_VSS_c_7_p N_CKN_c_268_n 5.38016e-19
cc_78 N_VSS_c_29_p N_CKN_c_272_n 2.21217e-19
cc_79 N_VSS_c_52_p N_CKN_c_272_n 0.00111539f
cc_80 N_VSS_c_3_p N_CKN_c_274_n 0.00220607f
cc_81 N_VSS_c_32_p N_CKN_c_274_n 8.60018e-19
cc_82 N_VSS_c_23_p N_CKN_c_274_n 2.36534e-19
cc_83 N_VSS_c_33_p N_CKN_c_274_n 7.62758e-19
cc_84 N_VSS_c_7_p N_CKN_c_274_n 0.00158805f
cc_85 N_VSS_c_85_p N_CKN_c_274_n 8.14378e-19
cc_86 N_VSS_c_38_p N_CKN_c_274_n 9.16986e-19
cc_87 N_VSS_c_29_p N_CKN_c_274_n 0.00110784f
cc_88 N_VSS_c_4_p N_D_XI5.X0_CG 0.00265616f
cc_89 N_VSS_c_89_p N_D_c_305_n 9.49637e-19
cc_90 N_VSS_XI5.X0_PGD N_D_c_306_n 3.8966e-19
cc_91 N_VSS_XI0.X0_PGD N_D_c_306_n 2.22031e-19
cc_92 N_VSS_c_3_p N_D_c_308_n 6.13924e-19
cc_93 N_VSS_c_23_p N_D_c_308_n 5.5494e-19
cc_94 N_VSS_c_20_p N_D_c_308_n 3.48267e-19
cc_95 N_VSS_c_4_p N_D_c_308_n 4.56568e-19
cc_96 N_VSS_c_3_p N_D_c_312_n 3.48267e-19
cc_97 N_VSS_c_23_p N_D_c_312_n 4.56568e-19
cc_98 N_VSS_c_20_p N_D_c_312_n 6.88619e-19
cc_99 N_VSS_c_4_p N_D_c_312_n 6.1245e-19
cc_100 N_VSS_XI4.X0_S N_X_XI5.X0_D 3.43419e-19
cc_101 N_VSS_c_45_p N_X_XI5.X0_D 3.48267e-19
cc_102 N_VSS_c_34_p N_X_XI0.X0_CG 0.00105235f
cc_103 N_VSS_XI5.X0_PGD N_X_c_334_n 2.09879e-19
cc_104 N_VSS_XI0.X0_PGD N_X_c_334_n 3.99472e-19
cc_105 N_VSS_c_38_p N_X_c_336_n 2.5064e-19
cc_106 N_VSS_XI4.X0_S N_X_c_337_n 3.48267e-19
cc_107 N_VSS_c_3_p N_X_c_337_n 4.71026e-19
cc_108 N_VSS_c_45_p N_X_c_337_n 5.69026e-19
cc_109 N_VSS_c_52_p N_X_c_337_n 2.04792e-19
cc_110 N_VSS_c_3_p N_X_c_341_n 0.00157847f
cc_111 N_VSS_c_52_p N_X_c_341_n 3.24972e-19
cc_112 N_VSS_c_3_p N_X_c_343_n 3.48267e-19
cc_113 N_VSS_c_4_p N_X_c_343_n 2.00604e-19
cc_114 N_VSS_XI3.X0_S N_Q_XI3.X0_D 3.43419e-19
cc_115 N_VSS_c_32_p N_Q_XI3.X0_D 3.48267e-19
cc_116 N_VSS_XI3.X0_S Q 3.48267e-19
cc_117 N_VSS_c_32_p Q 4.99861e-19
cc_118 N_CK_c_122_n N_VDD_XI1.X0_PGD 4.16623e-19
cc_119 N_CK_XI5.X0_PGS N_VDD_XI4.X0_PGD 2.40707e-19
cc_120 N_CK_c_123_n N_VDD_c_154_n 2.40707e-19
cc_121 CK N_VDD_c_155_n 5.04211e-19
cc_122 N_CK_c_129_p N_VDD_c_155_n 5.23418e-19
cc_123 N_CK_c_122_n N_VDD_c_159_n 0.00141086f
cc_124 CK N_VDD_c_159_n 0.00141439f
cc_125 N_CK_c_129_p N_VDD_c_159_n 0.00120361f
cc_126 N_CK_XI5.X0_PGS N_VDD_c_164_n 2.38687e-19
cc_127 N_CK_c_123_n N_VDD_c_164_n 5.38952e-19
cc_128 CK N_VDD_c_164_n 3.91916e-19
cc_129 N_CK_c_129_p N_VDD_c_164_n 2.80271e-19
cc_130 CK N_VDD_c_199_n 6.07878e-19
cc_131 N_CK_c_129_p N_VDD_c_199_n 4.67029e-19
cc_132 CK N_VDD_c_206_n 4.56568e-19
cc_133 N_CK_c_129_p N_VDD_c_206_n 0.00211811f
cc_134 N_CK_XI5.X0_PGS N_CKN_XI4.X0_PGS 4.11563e-19
cc_135 N_CK_XI5.X0_PGS N_CKN_c_283_n 2.73384e-19
cc_136 N_CK_XI5.X0_PGS N_D_XI5.X0_CG 4.28946e-19
cc_137 N_CK_XI5.X0_PGS N_D_XI4.X0_CG 2.59344e-19
cc_138 N_CK_XI5.X0_PGS N_D_c_312_n 0.00300565f
cc_139 N_CK_XI5.X0_PGS N_X_XI0.X0_CG 2.6404e-19
cc_140 N_CK_XI5.X0_PGS N_X_c_346_n 4.97357e-19
cc_141 N_CK_XI5.X0_PGS N_X_c_343_n 0.00630896f
cc_142 N_VDD_XI2.X0_S N_CKN_XI1.X0_D 3.43419e-19
cc_143 N_VDD_c_190_n N_CKN_XI4.X0_PGS 5.54393e-19
cc_144 N_VDD_c_190_n N_CKN_c_283_n 8.21431e-19
cc_145 N_VDD_XI2.X0_S N_CKN_c_268_n 3.48267e-19
cc_146 N_VDD_c_159_n N_CKN_c_268_n 5.01863e-19
cc_147 N_VDD_c_164_n N_CKN_c_268_n 5.35331e-19
cc_148 N_VDD_c_199_n N_CKN_c_268_n 6.42405e-19
cc_149 N_VDD_c_190_n N_CKN_c_272_n 7.71262e-19
cc_150 N_VDD_c_159_n N_CKN_c_274_n 4.68667e-19
cc_151 N_VDD_c_166_n N_CKN_c_274_n 3.15582e-19
cc_152 N_VDD_c_176_n N_CKN_c_274_n 4.71809e-19
cc_153 N_VDD_c_183_n N_CKN_c_274_n 2.56401e-19
cc_154 N_VDD_c_211_n N_D_XI4.X0_CG 0.00105644f
cc_155 N_VDD_XI3.X0_PGD N_D_c_306_n 2.08865e-19
cc_156 N_VDD_XI4.X0_PGD N_D_c_306_n 4.04053e-19
cc_157 N_VDD_XI2.X0_S N_X_XI5.X0_D 3.43419e-19
cc_158 N_VDD_c_164_n N_X_XI5.X0_D 3.48267e-19
cc_159 N_VDD_c_166_n N_X_XI5.X0_D 3.7884e-19
cc_160 N_VDD_c_208_n N_X_c_346_n 0.00269538f
cc_161 N_VDD_XI3.X0_PGD N_X_c_334_n 3.93054e-19
cc_162 N_VDD_XI4.X0_PGD N_X_c_334_n 2.22031e-19
cc_163 N_VDD_c_250_p N_X_c_354_n 8.95961e-19
cc_164 N_VDD_c_208_n N_X_c_354_n 2.97161e-19
cc_165 N_VDD_XI2.X0_S N_X_c_337_n 3.48267e-19
cc_166 N_VDD_c_164_n N_X_c_337_n 6.883e-19
cc_167 N_VDD_c_166_n N_X_c_337_n 5.3319e-19
cc_168 N_VDD_c_190_n N_X_c_337_n 8.74231e-19
cc_169 N_VDD_c_172_n N_X_c_341_n 6.5515e-19
cc_170 N_VDD_c_208_n N_X_c_341_n 4.80549e-19
cc_171 N_VDD_c_172_n N_X_c_343_n 4.85469e-19
cc_172 N_VDD_c_208_n N_X_c_343_n 6.1245e-19
cc_173 N_VDD_XI0.X0_S N_Q_XI3.X0_D 3.43419e-19
cc_174 N_VDD_c_176_n N_Q_XI3.X0_D 3.7884e-19
cc_175 N_VDD_c_188_n N_Q_XI3.X0_D 3.72199e-19
cc_176 N_VDD_XI0.X0_S Q 3.48267e-19
cc_177 N_VDD_c_176_n Q 5.12447e-19
cc_178 N_VDD_c_188_n Q 7.06537e-19
cc_179 N_CKN_XI4.X0_PGS N_D_XI4.X0_CG 0.00392964f
cc_180 N_CKN_XI4.X0_PGS N_X_c_334_n 0.00402435f
cc_181 N_CKN_c_283_n N_X_c_336_n 5.71169e-19
cc_182 N_CKN_c_274_n N_X_c_336_n 0.00120349f
cc_183 N_CKN_c_268_n N_X_c_337_n 2.66307e-19
cc_184 N_CKN_c_272_n N_X_c_337_n 8.08281e-19
cc_185 N_CKN_c_274_n N_X_c_337_n 6.2695e-19
cc_186 N_CKN_c_274_n N_X_c_341_n 7.98434e-19
cc_187 N_D_c_306_n N_X_c_334_n 0.00454934f
cc_188 N_D_c_306_n N_X_c_337_n 2.96904e-19
cc_189 N_D_c_308_n N_X_c_337_n 0.00151915f
cc_190 N_D_c_312_n N_X_c_337_n 9.22925e-19
cc_191 N_D_c_308_n N_X_c_341_n 0.00146206f
cc_192 N_D_c_312_n N_X_c_341_n 0.00103457f
cc_193 N_D_c_308_n N_X_c_343_n 4.56568e-19
cc_194 N_D_c_312_n N_X_c_343_n 0.00373298f
cc_195 N_X_c_336_n N_Q_XI3.X0_D 5.75967e-19
cc_196 N_X_c_336_n Q 8.57825e-19
*
.ends
*
*
.subckt DFFQ1_HPNW4 CK D Q VDD VSS
xgate (VSS CK VDD D Q) G3_DFFQ1_N1
.ends
*
* File: G1_INV1_N1.pex.netlist
* Created: Fri Feb 18 12:29:10 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G1_INV1_N1_VDD 2 5 15 28 30 34 37 43 Vss
c23 43 Vss 0.00628299f
c24 34 Vss 7.87399e-19
c25 30 Vss 0.00507852f
c26 28 Vss 0.00249774f
c27 26 Vss 0.00167323f
c28 15 Vss 0.0355813f
c29 14 Vss 0.102384f
c30 5 Vss 0.164813f
c31 2 Vss 0.00212755f
r32 34 43 1.16709
r33 32 34 2.45904
r34 31 37 0.326018
r35 30 32 0.652036
r36 30 31 7.41879
r37 26 37 0.326018
r38 26 28 5.08479
r39 17 43 0.214393
r40 15 17 1.4004
r41 14 18 0.652036
r42 14 17 1.5171
r43 11 15 0.652036
r44 5 18 2.5674
r45 5 11 2.5674
r46 2 28 1.16709
.ends

.subckt PM_G1_INV1_N1_A 2 4 9 12 22 25 28 Vss
c8 28 Vss 0.00718398f
c9 12 Vss 0.227852f
c10 9 Vss 0.0715834f
c11 7 Vss 0.0247918f
c12 4 Vss 0.0847975f
r13 25 28 1.16709
r14 22 25 0.0530455
r15 15 28 0.0476429
r16 13 15 0.326018
r17 13 15 0.1167
r18 12 16 0.652036
r19 12 15 6.7686
r20 9 28 0.357321
r21 7 15 0.326018
r22 7 9 0.40845
r23 4 16 2.5674
r24 2 9 2.15895
.ends

.subckt PM_G1_INV1_N1_VSS 3 6 14 27 32 37 49 50 56 Vss
c26 51 Vss 0.00126572f
c27 50 Vss 6.56738e-19
c28 49 Vss 0.00355297f
c29 37 Vss 0.0039192f
c30 32 Vss 0.00204286f
c31 27 Vss 6.63162e-19
c32 15 Vss 0.0358722f
c33 14 Vss 0.0994269f
c34 6 Vss 0.00276734f
c35 3 Vss 0.163777f
r36 51 56 0.326018
r37 49 56 0.326018
r38 49 50 7.46046
r39 45 50 0.652036
r40 32 51 5.08479
r41 27 37 1.16709
r42 27 45 2.41736
r43 17 37 0.238214
r44 15 17 1.45875
r45 14 18 0.652036
r46 14 17 1.45875
r47 11 15 0.652036
r48 6 32 1.16709
r49 3 18 2.5674
r50 3 11 2.5674
.ends

.subckt PM_G1_INV1_N1_Z 2 16 Vss
c11 2 Vss 0.00148239f
r12 16 19 0.125036
r13 2 19 1.16709
.ends

.subckt G1_INV1_N1  VDD A VSS Z
*
* Z	Z
* VSS	VSS
* A	A
* VDD	VDD
XI2.X0 N_Z_XI2.X0_D N_VSS_XI2.X0_PGD N_A_XI2.X0_CG N_VSS_XI2.X0_PGD
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI1.X0 N_Z_XI2.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW4
*
x_PM_G1_INV1_N1_VDD N_VDD_XI2.X0_S N_VDD_XI1.X0_PGD N_VDD_c_5_p N_VDD_c_4_p
+ N_VDD_c_6_p N_VDD_c_9_p VDD N_VDD_c_1_p Vss PM_G1_INV1_N1_VDD
x_PM_G1_INV1_N1_A N_A_XI2.X0_CG N_A_XI1.X0_CG N_A_c_29_p N_A_c_25_n A N_A_c_27_p
+ N_A_c_28_p Vss PM_G1_INV1_N1_A
x_PM_G1_INV1_N1_VSS N_VSS_XI2.X0_PGD N_VSS_XI1.X0_S N_VSS_c_34_n N_VSS_c_36_n
+ N_VSS_c_40_n N_VSS_c_42_n N_VSS_c_45_n N_VSS_c_46_n VSS Vss PM_G1_INV1_N1_VSS
x_PM_G1_INV1_N1_Z N_Z_XI2.X0_D Z Vss PM_G1_INV1_N1_Z
cc_1 N_VDD_c_1_p N_A_XI1.X0_CG 8.21222e-19
cc_2 N_VDD_XI1.X0_PGD N_A_c_25_n 4.26524e-19
cc_3 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00171093f
cc_4 N_VDD_c_4_p N_VSS_XI2.X0_PGD 4.197e-19
cc_5 N_VDD_c_5_p N_VSS_c_34_n 0.00171093f
cc_6 N_VDD_c_6_p N_VSS_c_34_n 4.82774e-19
cc_7 N_VDD_c_4_p N_VSS_c_36_n 0.00304634f
cc_8 N_VDD_c_6_p N_VSS_c_36_n 0.0015849f
cc_9 N_VDD_c_9_p N_VSS_c_36_n 9.51078e-19
cc_10 N_VDD_c_1_p N_VSS_c_36_n 3.5189e-19
cc_11 N_VDD_c_4_p N_VSS_c_40_n 3.08259e-19
cc_12 N_VDD_c_9_p N_VSS_c_40_n 0.00107037f
cc_13 N_VDD_c_4_p N_VSS_c_42_n 9.54992e-19
cc_14 N_VDD_c_9_p N_VSS_c_42_n 3.83199e-19
cc_15 N_VDD_c_1_p N_VSS_c_42_n 7.7548e-19
cc_16 N_VDD_c_6_p N_VSS_c_45_n 0.005791f
cc_17 N_VDD_c_6_p N_VSS_c_46_n 0.00172748f
cc_18 N_VDD_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_19 N_VDD_c_4_p N_Z_XI2.X0_D 3.48267e-19
cc_20 N_VDD_c_6_p N_Z_XI2.X0_D 3.55567e-19
cc_21 N_VDD_XI2.X0_S Z 3.48267e-19
cc_22 N_VDD_c_4_p Z 7.06424e-19
cc_23 N_VDD_c_6_p Z 4.789e-19
cc_24 N_A_c_25_n N_VSS_XI2.X0_PGD 4.21166e-19
cc_25 N_A_c_27_p N_VSS_c_36_n 0.00103813f
cc_26 N_A_c_28_p N_VSS_c_36_n 4.99367e-19
cc_27 N_A_c_29_p N_VSS_c_42_n 0.00250475f
cc_28 N_A_c_27_p N_VSS_c_42_n 4.99367e-19
cc_29 N_A_c_28_p N_VSS_c_42_n 0.0014909f
cc_30 N_VSS_XI1.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_31 N_VSS_c_40_n N_Z_XI2.X0_D 3.48267e-19
cc_32 N_VSS_XI1.X0_S Z 3.48267e-19
cc_33 N_VSS_c_40_n Z 7.85754e-19
cc_34 N_VSS_c_45_n Z 2.54816e-19
*
.ends
*
*
.subckt INV1_HPNW4 A Y VDD VSS
xgate (VDD A VSS Y) G1_INV1_N1
.ends
*
* File: G3_LATQ1_N1.pex.netlist
* Created: Tue Apr  5 11:43:13 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_LATQ1_N1_VDD 2 4 6 8 10 12 14 31 34 42 48 66 68 69 70 73 75 76 79
+ 81 85 89 91 92 94 100 105 Vss
c91 105 Vss 0.00462608f
c92 100 Vss 0.00538553f
c93 92 Vss 2.39889e-19
c94 91 Vss 3.56526e-19
c95 89 Vss 0.002537f
c96 87 Vss 0.00169593f
c97 85 Vss 9.25444e-19
c98 81 Vss 0.00432906f
c99 79 Vss 0.00113626f
c100 76 Vss 8.64506e-19
c101 75 Vss 0.00220359f
c102 73 Vss 0.00166444f
c103 70 Vss 8.63529e-19
c104 69 Vss 0.00558368f
c105 68 Vss 0.00685141f
c106 66 Vss 0.00204371f
c107 53 Vss 0.0307391f
c108 48 Vss 0.230209f
c109 42 Vss 0.0346914f
c110 41 Vss 0.0656875f
c111 34 Vss 6.95602e-20
c112 32 Vss 0.0348624f
c113 31 Vss 0.1003f
c114 14 Vss 0.0852073f
c115 12 Vss 0.00176834f
c116 10 Vss 0.0837105f
c117 8 Vss 0.0825478f
c118 6 Vss 0.0832227f
c119 4 Vss 0.0825437f
c120 2 Vss 0.00231819f
r121 87 94 0.326018
r122 87 89 4.83471
r123 85 105 1.16709
r124 83 85 2.16729
r125 82 92 0.494161
r126 81 94 0.326018
r127 81 82 7.41879
r128 79 100 1.16709
r129 77 92 0.128424
r130 77 79 2.16729
r131 75 92 0.494161
r132 75 76 4.41793
r133 71 91 0.0828784
r134 71 73 1.82344
r135 69 83 0.652036
r136 69 70 10.1279
r137 68 76 0.652036
r138 67 91 0.551426
r139 67 68 13.3371
r140 66 91 0.551426
r141 65 70 0.652036
r142 65 66 4.16786
r143 49 53 0.494161
r144 48 50 0.652036
r145 48 49 6.8853
r146 45 53 0.128424
r147 44 105 0.238214
r148 42 44 1.45875
r149 41 53 0.494161
r150 41 44 1.45875
r151 38 42 0.652036
r152 34 100 0.238214
r153 32 34 1.5171
r154 31 35 0.652036
r155 31 34 1.4004
r156 28 32 0.652036
r157 14 50 2.5674
r158 12 89 1.16709
r159 10 45 2.5674
r160 8 38 2.5674
r161 6 28 2.5674
r162 4 35 2.5674
r163 2 73 1.16709
.ends

.subckt PM_G3_LATQ1_N1_VSS 2 4 6 8 10 12 16 31 32 42 48 66 71 76 81 90 95 104
+ 106 107 108 113 114 119 129 130 132 Vss
c83 130 Vss 3.75522e-19
c84 129 Vss 4.28045e-19
c85 125 Vss 0.00127887f
c86 119 Vss 0.00326191f
c87 114 Vss 8.18866e-19
c88 113 Vss 0.00406272f
c89 108 Vss 8.24051e-19
c90 107 Vss 0.00164689f
c91 106 Vss 0.00145595f
c92 104 Vss 0.0042874f
c93 95 Vss 0.00390998f
c94 90 Vss 0.00430366f
c95 81 Vss 0.0025736f
c96 76 Vss 6.81193e-19
c97 71 Vss 9.80151e-19
c98 66 Vss 0.00132247f
c99 53 Vss 0.0307391f
c100 48 Vss 0.230436f
c101 42 Vss 0.0338877f
c102 41 Vss 0.0647949f
c103 32 Vss 0.0341879f
c104 31 Vss 0.0984533f
c105 16 Vss 0.085351f
c106 12 Vss 0.0838423f
c107 10 Vss 0.0825458f
c108 8 Vss 0.00178431f
c109 6 Vss 0.00237018f
c110 4 Vss 0.0842992f
c111 2 Vss 0.0825494f
r112 125 132 0.326018
r113 120 130 0.494161
r114 119 132 0.326018
r115 119 120 7.46046
r116 115 130 0.128424
r117 113 121 0.652036
r118 113 114 10.1279
r119 109 129 0.0828784
r120 107 130 0.494161
r121 107 108 4.37625
r122 106 114 0.652036
r123 105 129 0.551426
r124 105 106 4.16786
r125 104 129 0.551426
r126 103 108 0.652036
r127 103 104 13.3371
r128 81 125 4.83471
r129 76 95 1.16709
r130 76 121 2.16729
r131 71 90 1.16709
r132 71 115 2.16729
r133 66 109 1.82344
r134 49 53 0.494161
r135 48 50 0.652036
r136 48 49 6.8853
r137 45 53 0.128424
r138 44 95 0.238214
r139 42 44 1.45875
r140 41 53 0.494161
r141 41 44 1.45875
r142 38 42 0.652036
r143 34 90 0.238214
r144 32 34 1.45875
r145 31 35 0.652036
r146 31 34 1.45875
r147 28 32 0.652036
r148 16 50 2.5674
r149 12 45 2.5674
r150 10 38 2.5674
r151 8 81 1.16709
r152 6 66 1.16709
r153 4 28 2.5674
r154 2 35 2.5674
.ends

.subckt PM_G3_LATQ1_N1_G 2 4 6 14 15 22 31 37 Vss
c28 37 Vss 0.00243204f
c29 31 Vss 4.35685e-19
c30 29 Vss 0.0294543f
c31 22 Vss 0.152644f
c32 15 Vss 0.175771f
c33 14 Vss 3.53242e-19
c34 10 Vss 0.0247918f
c35 6 Vss 0.0835217f
c36 4 Vss 0.0840272f
c37 2 Vss 0.0715834f
r38 34 37 1.16709
r39 31 34 0.0833571
r40 23 29 0.494161
r41 22 24 0.652036
r42 22 23 4.84305
r43 19 29 0.128424
r44 18 37 0.0476429
r45 16 18 0.326018
r46 16 18 0.1167
r47 15 29 0.494161
r48 15 18 6.7686
r49 14 37 0.357321
r50 10 18 0.326018
r51 10 14 0.40845
r52 6 24 2.5674
r53 4 19 2.5674
r54 2 14 2.15895
.ends

.subckt PM_G3_LATQ1_N1_QN 2 4 6 8 17 20 23 40 45 48 53 69 Vss
c48 69 Vss 3.70906e-19
c49 53 Vss 0.0021144f
c50 48 Vss 0.00799496f
c51 45 Vss 0.00464908f
c52 40 Vss 7.75457e-19
c53 23 Vss 1.9003e-19
c54 20 Vss 0.213496f
c55 17 Vss 0.0714043f
c56 15 Vss 0.0247918f
c57 8 Vss 0.00402754f
c58 6 Vss 0.00402754f
c59 4 Vss 0.0829687f
r60 65 69 0.652036
r61 48 69 13.7956
r62 48 50 4.58464
r63 45 48 4.58464
r64 40 53 1.16709
r65 40 65 1.83386
r66 23 53 0.0476429
r67 21 23 0.326018
r68 21 23 0.1167
r69 20 24 0.652036
r70 20 23 6.7686
r71 17 53 0.357321
r72 15 23 0.326018
r73 15 17 0.40845
r74 8 50 1.16709
r75 6 45 1.16709
r76 4 24 2.5674
r77 2 17 2.15895
.ends

.subckt PM_G3_LATQ1_N1_GN 2 6 12 27 29 30 32 39 Vss
c46 39 Vss 0.00259221f
c47 32 Vss 2.5038e-19
c48 30 Vss 7.22041e-19
c49 29 Vss 0.00123575f
c50 27 Vss 9.12307e-19
c51 12 Vss 0.171268f
c52 6 Vss 0.17763f
c53 2 Vss 0.00172036f
r54 32 39 1.16709
r55 29 32 0.531835
r56 29 30 1.70882
r57 25 30 0.652036
r58 25 27 4.00114
r59 14 39 0.197068
r60 12 16 0.652036
r61 12 14 4.668
r62 6 16 5.835
r63 2 27 1.16709
.ends

.subckt PM_G3_LATQ1_N1_Q 2 18 Vss
c12 18 Vss 4.14768e-19
c13 2 Vss 0.00150258f
r14 2 18 1.16709
.ends

.subckt PM_G3_LATQ1_N1_D 2 4 10 14 Vss
c14 14 Vss 4.15825e-19
c15 10 Vss 1.35847e-19
c16 2 Vss 0.365962f
r17 14 17 0.0416786
r18 10 17 1.16709
r19 4 10 6.4185
r20 2 10 6.4185
.ends

.subckt G3_LATQ1_N1  VDD VSS G Q D
*
* D	D
* Q	Q
* G	G
* VSS	VSS
* VDD	VDD
XI2.X0 N_GN_XI2.X0_D N_VSS_XI2.X0_PGD N_G_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI0.X0 N_Q_XI0.X0_D N_VDD_XI0.X0_PGD N_QN_XI0.X0_CG N_VDD_XI0.X0_PGS
+ N_VSS_XI0.X0_S TIGFET_HPNW4
XI1.X0 N_GN_XI2.X0_D N_VDD_XI1.X0_PGD N_G_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI3.X0 N_Q_XI0.X0_D N_VSS_XI3.X0_PGD N_QN_XI3.X0_CG N_VSS_XI3.X0_PGS
+ N_VDD_XI3.X0_S TIGFET_HPNW4
XI5.X0 N_QN_XI5.X0_D N_VDD_XI5.X0_PGD N_D_XI5.X0_CG N_G_XI5.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI4.X0 N_QN_XI4.X0_D N_VSS_XI4.X0_PGD N_D_XI4.X0_CG N_GN_XI4.X0_PGS
+ N_VDD_XI3.X0_S TIGFET_HPNW4
*
x_PM_G3_LATQ1_N1_VDD N_VDD_XI2.X0_S N_VDD_XI0.X0_PGD N_VDD_XI0.X0_PGS
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI3.X0_S N_VDD_XI5.X0_PGD N_VDD_c_10_p
+ N_VDD_c_58_p N_VDD_c_7_p N_VDD_c_47_p N_VDD_c_16_p N_VDD_c_3_p N_VDD_c_8_p
+ N_VDD_c_38_p N_VDD_c_14_p N_VDD_c_15_p N_VDD_c_42_p N_VDD_c_20_p N_VDD_c_11_p
+ N_VDD_c_18_p N_VDD_c_5_p N_VDD_c_35_p N_VDD_c_41_p VDD N_VDD_c_23_p
+ N_VDD_c_19_p Vss PM_G3_LATQ1_N1_VDD
x_PM_G3_LATQ1_N1_VSS N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS N_VSS_XI0.X0_S
+ N_VSS_XI1.X0_S N_VSS_XI3.X0_PGD N_VSS_XI3.X0_PGS N_VSS_XI4.X0_PGD N_VSS_c_98_n
+ N_VSS_c_100_n N_VSS_c_101_n N_VSS_c_103_n N_VSS_c_104_n N_VSS_c_107_n
+ N_VSS_c_111_n N_VSS_c_115_n N_VSS_c_116_n N_VSS_c_120_n N_VSS_c_124_n
+ N_VSS_c_127_n N_VSS_c_128_n N_VSS_c_129_n N_VSS_c_130_n N_VSS_c_133_n
+ N_VSS_c_134_n N_VSS_c_135_n N_VSS_c_136_n VSS Vss PM_G3_LATQ1_N1_VSS
x_PM_G3_LATQ1_N1_G N_G_XI2.X0_CG N_G_XI1.X0_CG N_G_XI5.X0_PGS N_G_c_183_n
+ N_G_c_177_n N_G_c_179_n G N_G_c_181_n Vss PM_G3_LATQ1_N1_G
x_PM_G3_LATQ1_N1_QN N_QN_XI0.X0_CG N_QN_XI3.X0_CG N_QN_XI5.X0_D N_QN_XI4.X0_D
+ N_QN_c_205_n N_QN_c_206_n N_QN_c_208_n N_QN_c_210_n N_QN_c_213_n N_QN_c_215_n
+ N_QN_c_218_n N_QN_c_221_n Vss PM_G3_LATQ1_N1_QN
x_PM_G3_LATQ1_N1_GN N_GN_XI2.X0_D N_GN_XI4.X0_PGS N_GN_c_254_n N_GN_c_256_n
+ N_GN_c_279_n N_GN_c_285_n N_GN_c_260_n N_GN_c_262_n Vss PM_G3_LATQ1_N1_GN
x_PM_G3_LATQ1_N1_Q N_Q_XI0.X0_D Q Vss PM_G3_LATQ1_N1_Q
x_PM_G3_LATQ1_N1_D N_D_XI5.X0_CG N_D_XI4.X0_CG N_D_c_314_n D Vss
+ PM_G3_LATQ1_N1_D
cc_1 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.00175469f
cc_2 N_VDD_XI0.X0_PGS N_VSS_XI2.X0_PGS 2.27468e-19
cc_3 N_VDD_c_3_p N_VSS_XI0.X0_S 9.5668e-19
cc_4 N_VDD_XI0.X0_PGD N_VSS_XI3.X0_PGD 0.00173629f
cc_5 N_VDD_c_5_p N_VSS_XI3.X0_PGS 2.46127e-19
cc_6 N_VDD_XI5.X0_PGD N_VSS_XI4.X0_PGD 2.27468e-19
cc_7 N_VDD_c_7_p N_VSS_c_98_n 0.00175469f
cc_8 N_VDD_c_8_p N_VSS_c_98_n 3.60588e-19
cc_9 N_VDD_c_8_p N_VSS_c_100_n 3.60588e-19
cc_10 N_VDD_c_10_p N_VSS_c_101_n 0.00173629f
cc_11 N_VDD_c_11_p N_VSS_c_101_n 2.60334e-19
cc_12 N_VDD_c_5_p N_VSS_c_103_n 7.75484e-19
cc_13 N_VDD_c_3_p N_VSS_c_104_n 0.00165395f
cc_14 N_VDD_c_14_p N_VSS_c_104_n 7.6714e-19
cc_15 N_VDD_c_15_p N_VSS_c_104_n 5.16845e-19
cc_16 N_VDD_c_16_p N_VSS_c_107_n 4.43871e-19
cc_17 N_VDD_c_8_p N_VSS_c_107_n 0.00161703f
cc_18 N_VDD_c_18_p N_VSS_c_107_n 9.31718e-19
cc_19 N_VDD_c_19_p N_VSS_c_107_n 3.48267e-19
cc_20 N_VDD_c_20_p N_VSS_c_111_n 9.36729e-19
cc_21 N_VDD_c_11_p N_VSS_c_111_n 0.00141228f
cc_22 N_VDD_c_5_p N_VSS_c_111_n 0.00291977f
cc_23 N_VDD_c_23_p N_VSS_c_111_n 3.5189e-19
cc_24 N_VDD_c_18_p N_VSS_c_115_n 0.00102583f
cc_25 N_VDD_c_16_p N_VSS_c_116_n 3.66936e-19
cc_26 N_VDD_c_8_p N_VSS_c_116_n 2.03837e-19
cc_27 N_VDD_c_18_p N_VSS_c_116_n 3.99794e-19
cc_28 N_VDD_c_19_p N_VSS_c_116_n 8.07896e-19
cc_29 N_VDD_c_20_p N_VSS_c_120_n 3.86045e-19
cc_30 N_VDD_c_11_p N_VSS_c_120_n 0.00112249f
cc_31 N_VDD_c_5_p N_VSS_c_120_n 9.54992e-19
cc_32 N_VDD_c_23_p N_VSS_c_120_n 8.1718e-19
cc_33 N_VDD_c_16_p N_VSS_c_124_n 0.00303537f
cc_34 N_VDD_c_3_p N_VSS_c_124_n 0.00544275f
cc_35 N_VDD_c_35_p N_VSS_c_124_n 0.00116512f
cc_36 N_VDD_c_3_p N_VSS_c_127_n 0.00305967f
cc_37 N_VDD_c_8_p N_VSS_c_128_n 0.00343927f
cc_38 N_VDD_c_38_p N_VSS_c_129_n 0.00106317f
cc_39 N_VDD_c_15_p N_VSS_c_130_n 0.00355199f
cc_40 N_VDD_c_11_p N_VSS_c_130_n 0.00567045f
cc_41 N_VDD_c_41_p N_VSS_c_130_n 9.48532e-19
cc_42 N_VDD_c_42_p N_VSS_c_133_n 0.00105938f
cc_43 N_VDD_c_8_p N_VSS_c_134_n 0.00557463f
cc_44 N_VDD_c_3_p N_VSS_c_135_n 8.91588e-19
cc_45 N_VDD_c_8_p N_VSS_c_136_n 7.74609e-19
cc_46 N_VDD_c_19_p N_G_XI1.X0_CG 8.09841e-19
cc_47 N_VDD_c_47_p N_G_XI5.X0_PGS 0.00162079f
cc_48 N_VDD_XI0.X0_PGD N_G_c_177_n 2.22031e-19
cc_49 N_VDD_XI1.X0_PGD N_G_c_177_n 3.93641e-19
cc_50 N_VDD_XI1.X0_PGS N_G_c_179_n 4.05198e-19
cc_51 N_VDD_c_3_p G 3.46645e-19
cc_52 N_VDD_c_3_p N_G_c_181_n 4.43544e-19
cc_53 N_VDD_XI3.X0_S N_QN_XI4.X0_D 3.43419e-19
cc_54 N_VDD_c_5_p N_QN_XI4.X0_D 3.48267e-19
cc_55 N_VDD_c_23_p N_QN_c_205_n 0.00269246f
cc_56 N_VDD_XI0.X0_PGD N_QN_c_206_n 4.05198e-19
cc_57 N_VDD_XI1.X0_PGD N_QN_c_206_n 2.0936e-19
cc_58 N_VDD_c_58_p N_QN_c_208_n 9.69462e-19
cc_59 N_VDD_c_23_p N_QN_c_208_n 2.60536e-19
cc_60 N_VDD_c_3_p N_QN_c_210_n 4.49462e-19
cc_61 N_VDD_c_20_p N_QN_c_210_n 4.57093e-19
cc_62 N_VDD_c_23_p N_QN_c_210_n 4.4444e-19
cc_63 N_VDD_XI3.X0_S N_QN_c_213_n 3.48267e-19
cc_64 N_VDD_c_5_p N_QN_c_213_n 9.00822e-19
cc_65 N_VDD_c_8_p N_QN_c_215_n 4.48879e-19
cc_66 N_VDD_c_11_p N_QN_c_215_n 3.93728e-19
cc_67 N_VDD_c_5_p N_QN_c_215_n 3.58217e-19
cc_68 N_VDD_c_3_p N_QN_c_218_n 6.61926e-19
cc_69 N_VDD_c_20_p N_QN_c_218_n 4.85469e-19
cc_70 N_VDD_c_23_p N_QN_c_218_n 6.1245e-19
cc_71 N_VDD_c_3_p N_QN_c_221_n 4.64547e-19
cc_72 N_VDD_XI2.X0_S N_GN_XI2.X0_D 3.43419e-19
cc_73 N_VDD_c_8_p N_GN_XI2.X0_D 3.7884e-19
cc_74 N_VDD_c_14_p N_GN_XI2.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_PGS N_GN_c_254_n 3.40151e-19
cc_76 N_VDD_c_47_p N_GN_c_254_n 3.20239e-19
cc_77 N_VDD_XI2.X0_S N_GN_c_256_n 3.48267e-19
cc_78 N_VDD_c_3_p N_GN_c_256_n 6.12365e-19
cc_79 N_VDD_c_8_p N_GN_c_256_n 5.32769e-19
cc_80 N_VDD_c_14_p N_GN_c_256_n 7.89245e-19
cc_81 N_VDD_c_18_p N_GN_c_260_n 2.2082e-19
cc_82 N_VDD_c_19_p N_GN_c_260_n 2.46105e-19
cc_83 N_VDD_c_18_p N_GN_c_262_n 2.68489e-19
cc_84 N_VDD_c_19_p N_GN_c_262_n 5.71759e-19
cc_85 N_VDD_XI3.X0_S N_Q_XI0.X0_D 3.43419e-19
cc_86 N_VDD_c_11_p N_Q_XI0.X0_D 3.7884e-19
cc_87 N_VDD_c_5_p N_Q_XI0.X0_D 3.48267e-19
cc_88 N_VDD_XI3.X0_S Q 3.48267e-19
cc_89 N_VDD_c_11_p Q 5.12447e-19
cc_90 N_VDD_c_5_p Q 7.06424e-19
cc_91 N_VDD_c_47_p N_D_XI5.X0_CG 4.07085e-19
cc_92 N_VSS_c_116_n N_G_XI2.X0_CG 0.00265616f
cc_93 N_VSS_c_116_n N_G_c_183_n 9.49637e-19
cc_94 N_VSS_XI2.X0_PGD N_G_c_177_n 3.99472e-19
cc_95 N_VSS_XI3.X0_PGD N_G_c_177_n 2.0936e-19
cc_96 N_VSS_c_107_n G 5.5494e-19
cc_97 N_VSS_c_116_n G 4.56568e-19
cc_98 N_VSS_c_124_n G 3.38887e-19
cc_99 N_VSS_c_107_n N_G_c_181_n 4.56568e-19
cc_100 N_VSS_c_116_n N_G_c_181_n 6.1245e-19
cc_101 N_VSS_c_120_n N_QN_XI3.X0_CG 8.05748e-19
cc_102 N_VSS_XI1.X0_S N_QN_XI5.X0_D 3.43419e-19
cc_103 N_VSS_c_115_n N_QN_XI5.X0_D 3.48267e-19
cc_104 N_VSS_XI2.X0_PGD N_QN_c_206_n 2.22031e-19
cc_105 N_VSS_XI3.X0_PGD N_QN_c_206_n 3.89061e-19
cc_106 N_VSS_c_130_n N_QN_c_210_n 2.91026e-19
cc_107 N_VSS_c_115_n N_QN_c_213_n 8.97415e-19
cc_108 N_VSS_c_111_n N_QN_c_215_n 3.5258e-19
cc_109 N_VSS_c_115_n N_QN_c_215_n 7.99552e-19
cc_110 N_VSS_c_130_n N_QN_c_215_n 6.85871e-19
cc_111 N_VSS_c_134_n N_QN_c_215_n 9.55516e-19
cc_112 N_VSS_c_107_n N_QN_c_221_n 5.43247e-19
cc_113 N_VSS_c_124_n N_QN_c_221_n 0.00168288f
cc_114 N_VSS_XI1.X0_S N_GN_XI2.X0_D 3.43419e-19
cc_115 N_VSS_c_115_n N_GN_XI2.X0_D 3.48267e-19
cc_116 N_VSS_c_103_n N_GN_XI4.X0_PGS 0.00163489f
cc_117 N_VSS_XI3.X0_PGS N_GN_c_254_n 6.77138e-19
cc_118 N_VSS_c_103_n N_GN_c_254_n 2.57527e-19
cc_119 N_VSS_XI1.X0_S N_GN_c_256_n 3.48267e-19
cc_120 N_VSS_c_115_n N_GN_c_256_n 4.97497e-19
cc_121 N_VSS_c_124_n N_GN_c_256_n 4.46497e-19
cc_122 N_VSS_c_120_n N_GN_c_260_n 2.46105e-19
cc_123 N_VSS_c_111_n N_GN_c_262_n 2.52506e-19
cc_124 N_VSS_c_120_n N_GN_c_262_n 5.99566e-19
cc_125 N_VSS_XI0.X0_S N_Q_XI0.X0_D 3.43419e-19
cc_126 N_VSS_c_104_n N_Q_XI0.X0_D 3.48267e-19
cc_127 N_VSS_XI0.X0_S Q 3.48267e-19
cc_128 N_VSS_c_104_n Q 7.78122e-19
cc_129 N_VSS_c_103_n N_D_XI5.X0_CG 4.07085e-19
cc_130 N_G_c_177_n N_QN_c_206_n 0.003965f
cc_131 G N_QN_c_210_n 5.07332e-19
cc_132 N_G_c_181_n N_QN_c_210_n 4.54925e-19
cc_133 N_G_c_181_n N_QN_c_218_n 0.00269321f
cc_134 N_G_c_179_n N_GN_c_254_n 0.00851239f
cc_135 N_G_c_177_n N_GN_c_256_n 3.2445e-19
cc_136 G N_GN_c_256_n 0.00153131f
cc_137 N_G_c_181_n N_GN_c_256_n 9.18093e-19
cc_138 N_G_c_177_n N_GN_c_279_n 3.7133e-19
cc_139 N_G_c_177_n N_GN_c_262_n 9.94034e-19
cc_140 N_G_c_181_n N_GN_c_262_n 2.41671e-19
cc_141 N_G_XI5.X0_PGS N_D_XI5.X0_CG 0.00409312f
cc_142 N_QN_c_206_n N_GN_XI4.X0_PGS 0.00182388f
cc_143 N_QN_c_213_n N_GN_c_256_n 7.80248e-19
cc_144 N_QN_c_215_n N_GN_c_279_n 8.96813e-19
cc_145 N_QN_c_215_n N_GN_c_285_n 0.00118168f
cc_146 N_QN_c_215_n N_GN_c_260_n 9.24681e-19
cc_147 N_QN_c_206_n N_GN_c_262_n 8.57779e-19
cc_148 N_QN_c_218_n N_GN_c_262_n 2.75519e-19
cc_149 N_QN_c_206_n N_D_XI5.X0_CG 3.26559e-19
cc_150 N_QN_c_213_n N_D_XI5.X0_CG 0.00101289f
cc_151 N_QN_c_213_n N_D_c_314_n 0.00127983f
cc_152 N_QN_c_213_n D 0.00141415f
cc_153 N_QN_c_215_n D 0.00146947f
cc_154 N_GN_c_285_n N_Q_XI0.X0_D 5.19956e-19
cc_155 N_GN_c_285_n Q 6.79271e-19
cc_156 N_GN_XI4.X0_PGS N_D_XI5.X0_CG 0.00503657f
cc_157 N_GN_c_254_n N_D_c_314_n 0.00333193f
cc_158 N_GN_c_260_n N_D_c_314_n 3.73302e-19
cc_159 N_GN_c_262_n N_D_c_314_n 8.5422e-19
cc_160 N_GN_c_260_n D 2.88184e-19
cc_161 N_GN_c_262_n D 3.48267e-19
*
.ends
*
*
.subckt LATQ1_HPNW4 D G Q VDD VSS
xgate (VDD VSS G Q D) G3_LATQ1_N1
.ends
*
* File: G4_MAJ3_N1.pex.netlist
* Created: Wed Mar  2 17:07:12 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MAJ3_N1_VDD 2 4 7 11 27 28 31 32 51 52 54 56 57 61 65 67 68 71 75
+ 78 79 80 90 95 Vss
c80 95 Vss 0.00471931f
c81 90 Vss 0.00455939f
c82 80 Vss 3.56526e-19
c83 79 Vss 3.56526e-19
c84 75 Vss 3.84406e-19
c85 71 Vss 9.33011e-19
c86 68 Vss 8.63529e-19
c87 67 Vss 0.00539264f
c88 65 Vss 0.00133146f
c89 61 Vss 0.00133512f
c90 57 Vss 0.00563423f
c91 56 Vss 0.0019972f
c92 54 Vss 0.00437281f
c93 52 Vss 0.00204371f
c94 51 Vss 8.63529e-19
c95 32 Vss 0.0336444f
c96 31 Vss 0.0988545f
c97 28 Vss 0.0346129f
c98 27 Vss 0.0990038f
c99 11 Vss 0.165071f
c100 7 Vss 0.165416f
c101 4 Vss 0.00207958f
c102 2 Vss 0.0026194f
r103 75 95 1.16709
r104 73 75 2.16729
r105 71 90 1.16709
r106 69 71 2.16729
r107 67 73 0.652036
r108 67 68 10.1279
r109 63 80 0.0828784
r110 63 65 1.82344
r111 59 79 0.0828784
r112 59 61 1.82344
r113 58 78 0.326018
r114 57 69 0.652036
r115 57 58 10.1279
r116 56 68 0.652036
r117 55 80 0.551426
r118 55 56 4.16786
r119 54 80 0.551426
r120 53 79 0.551426
r121 53 54 7.83557
r122 52 79 0.551426
r123 51 78 0.326018
r124 51 52 4.16786
r125 34 95 0.238214
r126 32 34 1.45875
r127 31 38 0.652036
r128 31 34 1.45875
r129 30 90 0.238214
r130 28 30 1.45875
r131 27 35 0.652036
r132 27 30 1.45875
r133 24 32 0.652036
r134 21 28 0.652036
r135 11 38 2.5674
r136 11 24 2.5674
r137 7 35 2.5674
r138 7 21 2.5674
r139 4 65 1.16709
r140 2 61 1.16709
.ends

.subckt PM_G4_MAJ3_N1_VSS 3 7 10 12 27 28 31 32 34 52 57 62 67 70 73 78 91 92 93
+ 94 95 104 114 115 117 Vss
c89 115 Vss 3.75522e-19
c90 114 Vss 3.75522e-19
c91 110 Vss 0.00127887f
c92 104 Vss 0.00344356f
c93 95 Vss 8.24051e-19
c94 94 Vss 0.00149351f
c95 93 Vss 8.24051e-19
c96 92 Vss 0.00149351f
c97 91 Vss 0.00617495f
c98 78 Vss 0.00390682f
c99 73 Vss 0.00498746f
c100 70 Vss 0.00347745f
c101 67 Vss 0.00294127f
c102 62 Vss 0.00184732f
c103 57 Vss 0.00132425f
c104 52 Vss 0.00115907f
c105 32 Vss 0.033157f
c106 31 Vss 0.0974849f
c107 28 Vss 0.0341879f
c108 27 Vss 0.0984533f
c109 12 Vss 0.00257143f
c110 10 Vss 0.00203161f
c111 7 Vss 0.166925f
c112 3 Vss 0.166819f
r113 110 117 0.326018
r114 106 115 0.494161
r115 105 114 0.494161
r116 104 117 0.326018
r117 104 105 7.46046
r118 100 115 0.128424
r119 96 114 0.128424
r120 94 115 0.494161
r121 94 95 4.37625
r122 92 114 0.494161
r123 92 93 4.37625
r124 91 95 0.652036
r125 90 93 0.652036
r126 90 91 18.8387
r127 70 106 8.04396
r128 67 70 5.41821
r129 62 110 4.83471
r130 57 78 1.16709
r131 57 100 2.16729
r132 52 73 1.16709
r133 52 96 2.16729
r134 34 78 0.238214
r135 32 34 1.45875
r136 31 38 0.652036
r137 31 34 1.45875
r138 30 73 0.238214
r139 28 30 1.45875
r140 27 35 0.652036
r141 27 30 1.45875
r142 24 32 0.652036
r143 21 28 0.652036
r144 12 67 1.16709
r145 10 62 1.16709
r146 7 38 2.5674
r147 7 24 2.5674
r148 3 35 2.5674
r149 3 21 2.5674
.ends

.subckt PM_G4_MAJ3_N1_A 2 4 6 8 11 15 29 32 53 57 69 72 74 77 79 81 82 85 87 90
+ 98 107 Vss
c80 110 Vss 1.14262e-19
c81 107 Vss 0.00533929f
c82 98 Vss 0.00481087f
c83 94 Vss 7.48717e-19
c84 87 Vss 6.11441e-19
c85 85 Vss 8.50217e-19
c86 82 Vss 4.65536e-19
c87 81 Vss 0.00274588f
c88 79 Vss 0.00488819f
c89 77 Vss 8.85587e-19
c90 74 Vss 0.00117147f
c91 73 Vss 0.00146569f
c92 72 Vss 0.00379017f
c93 69 Vss 0.00539132f
c94 57 Vss 0.135015f
c95 53 Vss 0.128028f
c96 32 Vss 0.2139f
c97 29 Vss 0.0749894f
c98 27 Vss 0.0247918f
c99 11 Vss 1.01176f
c100 8 Vss 0.00236553f
c101 6 Vss 0.00271742f
c102 4 Vss 0.0850321f
r103 107 110 0.1
r104 96 107 1.16709
r105 92 98 1.16709
r106 90 92 0.166714
r107 87 90 0.166714
r108 83 85 2.16729
r109 82 96 0.531835
r110 81 83 0.652036
r111 81 82 1.70882
r112 80 94 0.494161
r113 79 96 0.531835
r114 79 80 7.46046
r115 75 94 0.128424
r116 75 77 2.16729
r117 73 94 0.494161
r118 73 74 1.83386
r119 71 74 0.652036
r120 71 72 8.00229
r121 70 87 0.0685365
r122 69 72 0.652036
r123 69 70 10.2113
r124 55 57 4.53833
r125 52 110 0.262036
r126 52 53 2.26917
r127 49 52 2.26917
r128 44 57 0.00605528
r129 43 53 0.00605528
r130 40 55 0.00605528
r131 39 49 0.00605528
r132 35 98 0.0952857
r133 33 35 0.326018
r134 33 35 0.1167
r135 32 36 0.652036
r136 32 35 6.7686
r137 29 35 0.3335
r138 27 35 0.326018
r139 27 29 0.2334
r140 15 44 2.5674
r141 15 40 2.5674
r142 11 15 12.837
r143 11 43 2.5674
r144 11 15 12.837
r145 11 39 2.5674
r146 8 85 1.16709
r147 6 77 1.16709
r148 4 36 2.5674
r149 2 29 2.334
.ends

.subckt PM_G4_MAJ3_N1_BI 2 6 8 21 32 37 42 52 57 66 72 73 Vss
c61 73 Vss 3.33918e-19
c62 72 Vss 7.31231e-19
c63 66 Vss 0.00174781f
c64 57 Vss 0.00147766f
c65 52 Vss 0.00140496f
c66 42 Vss 0.0015273f
c67 37 Vss 0.00542097f
c68 32 Vss 0.00210957f
c69 21 Vss 0.0573997f
c70 6 Vss 0.0573997f
c71 2 Vss 0.0015046f
r72 72 73 0.65228
r73 71 72 3.42052
r74 66 71 0.65409
r75 42 57 1.16709
r76 42 73 2.1395
r77 37 52 1.16709
r78 37 77 12.0712
r79 37 66 1.96931
r80 32 49 1.16709
r81 32 77 2.08393
r82 21 57 0.50025
r83 18 52 0.50025
r84 8 21 1.80885
r85 6 18 1.80885
r86 2 49 0.1
.ends

.subckt PM_G4_MAJ3_N1_AI 2 7 11 31 37 46 51 60 69 Vss
c47 69 Vss 2.51637e-19
c48 60 Vss 0.00575758f
c49 51 Vss 0.00577434f
c50 46 Vss 9.64269e-19
c51 37 Vss 0.127837f
c52 36 Vss 1.23462e-19
c53 31 Vss 0.133405f
c54 7 Vss 1.0035f
c55 2 Vss 0.0015046f
r56 65 69 0.652036
r57 60 63 0.1
r58 51 63 1.16709
r59 51 69 13.7539
r60 46 65 2.16729
r61 36 60 0.262036
r62 36 37 2.334
r63 33 36 2.20433
r64 29 31 4.53833
r65 26 37 0.00605528
r66 25 31 0.00605528
r67 22 33 0.00605528
r68 21 29 0.00605528
r69 11 26 2.5674
r70 11 22 2.5674
r71 7 11 12.837
r72 7 25 2.5674
r73 7 11 12.837
r74 7 21 2.5674
r75 2 46 1.16709
.ends

.subckt PM_G4_MAJ3_N1_B 2 4 6 8 16 17 26 38 42 45 50 55 60 65 73 74 80 87 92 93
+ Vss
c73 93 Vss 4.59352e-19
c74 92 Vss 0.00214833f
c75 87 Vss 7.9499e-19
c76 80 Vss 8.69209e-19
c77 74 Vss 2.46868e-19
c78 73 Vss 0.00310209f
c79 65 Vss 0.00148695f
c80 60 Vss 0.00103393f
c81 55 Vss 0.004462f
c82 50 Vss 0.00190521f
c83 45 Vss 8.22554e-19
c84 38 Vss 0.00131454f
c85 26 Vss 0.0573997f
c86 20 Vss 0.0247918f
c87 17 Vss 0.0343999f
c88 16 Vss 0.183114f
c89 8 Vss 0.0573997f
c90 4 Vss 0.0714013f
c91 2 Vss 0.0847975f
r92 91 93 0.65228
r93 91 92 3.46076
r94 87 92 0.65228
r95 83 87 2.1006
r96 80 83 2.04225
r97 73 80 0.0685365
r98 73 74 10.3363
r99 69 74 0.652036
r100 50 65 1.16709
r101 50 93 2.1395
r102 45 60 1.16709
r103 45 83 0.0416786
r104 38 55 1.16709
r105 38 69 2.16729
r106 38 42 0.0833571
r107 36 55 0.0476429
r108 33 65 0.50025
r109 26 60 0.50025
r110 24 55 0.357321
r111 20 36 0.326018
r112 20 24 0.40845
r113 17 36 6.7686
r114 16 36 0.326018
r115 16 36 0.1167
r116 13 17 0.652036
r117 8 33 1.80885
r118 6 26 1.80885
r119 4 24 2.15895
r120 2 13 2.5674
.ends

.subckt PM_G4_MAJ3_N1_C 2 4 20 25 50 54 57 Vss
c27 57 Vss 0.00412628f
c28 54 Vss 7.72795e-19
c29 25 Vss 0.00139119f
c30 20 Vss 6.60907e-19
c31 4 Vss 0.00277614f
c32 2 Vss 0.00222834f
r33 50 57 1.08364
r34 50 54 9.25264
r35 25 57 0.521797
r36 20 54 0.521797
r37 4 25 1.16709
r38 2 20 1.16709
.ends

.subckt PM_G4_MAJ3_N1_Z 2 4 30 33 Vss
c33 30 Vss 0.00258707f
c34 4 Vss 0.00153036f
c35 2 Vss 0.00148239f
r36 33 35 4.50129
r37 30 33 4.668
r38 4 35 1.16709
r39 2 30 1.16709
.ends

.subckt G4_MAJ3_N1  VDD VSS A B C Z
*
* Z	Z
* C	C
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI6.X0 N_BI_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW4
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI5.X0 N_VSS_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_BI_XI6.X0_D TIGFET_HPNW4
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW4
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_BI_XI2.X0_CG N_AI_XI2.X0_PGD N_A_XI2.X0_S
+ TIGFET_HPNW4
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_B_XI4.X0_CG N_AI_XI4.X0_PGD N_C_XI4.X0_S
+ TIGFET_HPNW4
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_B_XI3.X0_CG N_A_XI3.X0_PGD N_A_XI3.X0_S
+ TIGFET_HPNW4
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_BI_XI1.X0_CG N_A_XI1.X0_PGD N_C_XI1.X0_S
+ TIGFET_HPNW4
*
x_PM_G4_MAJ3_N1_VDD N_VDD_XI6.X0_S N_VDD_XI8.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI7.X0_PGD N_VDD_c_65_p N_VDD_c_3_p N_VDD_c_66_p N_VDD_c_6_p
+ N_VDD_c_37_p N_VDD_c_9_p N_VDD_c_31_p N_VDD_c_13_p N_VDD_c_4_p N_VDD_c_36_p
+ N_VDD_c_38_p N_VDD_c_7_p N_VDD_c_40_p N_VDD_c_11_p N_VDD_c_15_p VDD
+ N_VDD_c_33_p N_VDD_c_34_p N_VDD_c_12_p N_VDD_c_16_p Vss PM_G4_MAJ3_N1_VDD
x_PM_G4_MAJ3_N1_VSS N_VSS_XI6.X0_PGD N_VSS_XI8.X0_PGD N_VSS_XI5.X0_D
+ N_VSS_XI7.X0_S N_VSS_c_83_n N_VSS_c_85_n N_VSS_c_86_n N_VSS_c_88_n
+ N_VSS_c_135_p N_VSS_c_89_n N_VSS_c_93_n N_VSS_c_97_n N_VSS_c_98_n
+ N_VSS_c_101_n N_VSS_c_102_n N_VSS_c_106_n N_VSS_c_110_n N_VSS_c_115_n
+ N_VSS_c_117_n N_VSS_c_118_n N_VSS_c_120_n N_VSS_c_121_n N_VSS_c_122_n
+ N_VSS_c_123_n VSS Vss PM_G4_MAJ3_N1_VSS
x_PM_G4_MAJ3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI2.X0_S N_A_XI3.X0_S
+ N_A_XI3.X0_PGD N_A_XI1.X0_PGD N_A_c_182_n N_A_c_171_n N_A_c_211_p N_A_c_213_p
+ N_A_c_172_n N_A_c_189_n N_A_c_177_n N_A_c_233_p N_A_c_199_p N_A_c_237_p
+ N_A_c_225_p N_A_c_236_p N_A_c_179_n A N_A_c_180_n N_A_c_207_p Vss
+ PM_G4_MAJ3_N1_A
x_PM_G4_MAJ3_N1_BI N_BI_XI6.X0_D N_BI_XI2.X0_CG N_BI_XI1.X0_CG N_BI_c_265_n
+ N_BI_c_253_n N_BI_c_262_n N_BI_c_269_n N_BI_c_270_n N_BI_c_271_n N_BI_c_273_n
+ N_BI_c_293_p N_BI_c_296_p Vss PM_G4_MAJ3_N1_BI
x_PM_G4_MAJ3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_315_n
+ N_AI_c_316_n N_AI_c_317_n N_AI_c_320_n N_AI_c_330_n N_AI_c_321_n Vss
+ PM_G4_MAJ3_N1_AI
x_PM_G4_MAJ3_N1_B N_B_XI6.X0_CG N_B_XI5.X0_CG N_B_XI4.X0_CG N_B_XI3.X0_CG
+ N_B_c_359_n N_B_c_377_n N_B_c_414_n N_B_c_361_n B N_B_c_380_n N_B_c_381_n
+ N_B_c_364_n N_B_c_386_n N_B_c_387_n N_B_c_371_n N_B_c_372_n N_B_c_405_n
+ N_B_c_408_n N_B_c_411_n N_B_c_412_n Vss PM_G4_MAJ3_N1_B
x_PM_G4_MAJ3_N1_C N_C_XI4.X0_S N_C_XI1.X0_S N_C_c_433_n N_C_c_435_n C
+ N_C_c_437_n N_C_c_436_n Vss PM_G4_MAJ3_N1_C
x_PM_G4_MAJ3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_463_n Z Vss PM_G4_MAJ3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017247f
cc_2 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172036f
cc_3 N_VDD_c_3_p N_VSS_c_83_n 0.0017247f
cc_4 N_VDD_c_4_p N_VSS_c_83_n 2.74208e-19
cc_5 N_VDD_c_4_p N_VSS_c_85_n 3.60588e-19
cc_6 N_VDD_c_6_p N_VSS_c_86_n 0.00172036f
cc_7 N_VDD_c_7_p N_VSS_c_86_n 2.46461e-19
cc_8 N_VDD_c_7_p N_VSS_c_88_n 3.60588e-19
cc_9 N_VDD_c_9_p N_VSS_c_89_n 4.43871e-19
cc_10 N_VDD_c_4_p N_VSS_c_89_n 0.00161703f
cc_11 N_VDD_c_11_p N_VSS_c_89_n 9.28314e-19
cc_12 N_VDD_c_12_p N_VSS_c_89_n 3.48267e-19
cc_13 N_VDD_c_13_p N_VSS_c_93_n 4.43871e-19
cc_14 N_VDD_c_7_p N_VSS_c_93_n 0.00161703f
cc_15 N_VDD_c_15_p N_VSS_c_93_n 8.31866e-19
cc_16 N_VDD_c_16_p N_VSS_c_93_n 3.48267e-19
cc_17 N_VDD_c_11_p N_VSS_c_97_n 8.49247e-19
cc_18 N_VDD_XI7.X0_PGD N_VSS_c_98_n 3.41313e-19
cc_19 N_VDD_c_15_p N_VSS_c_98_n 0.00507115f
cc_20 N_VDD_c_16_p N_VSS_c_98_n 9.58524e-19
cc_21 N_VDD_c_7_p N_VSS_c_101_n 0.00403287f
cc_22 N_VDD_c_9_p N_VSS_c_102_n 3.66936e-19
cc_23 N_VDD_c_4_p N_VSS_c_102_n 2.03837e-19
cc_24 N_VDD_c_11_p N_VSS_c_102_n 3.99794e-19
cc_25 N_VDD_c_12_p N_VSS_c_102_n 8.07896e-19
cc_26 N_VDD_c_13_p N_VSS_c_106_n 3.66936e-19
cc_27 N_VDD_c_7_p N_VSS_c_106_n 2.03837e-19
cc_28 N_VDD_c_15_p N_VSS_c_106_n 3.99794e-19
cc_29 N_VDD_c_16_p N_VSS_c_106_n 8.03027e-19
cc_30 N_VDD_c_9_p N_VSS_c_110_n 0.00303537f
cc_31 N_VDD_c_31_p N_VSS_c_110_n 0.00599011f
cc_32 N_VDD_c_13_p N_VSS_c_110_n 0.00284565f
cc_33 N_VDD_c_33_p N_VSS_c_110_n 0.00104624f
cc_34 N_VDD_c_34_p N_VSS_c_110_n 0.0010706f
cc_35 N_VDD_c_4_p N_VSS_c_115_n 0.00345066f
cc_36 N_VDD_c_36_p N_VSS_c_115_n 2.07484e-19
cc_37 N_VDD_c_37_p N_VSS_c_117_n 0.00106317f
cc_38 N_VDD_c_38_p N_VSS_c_118_n 2.07484e-19
cc_39 N_VDD_c_7_p N_VSS_c_118_n 0.00345066f
cc_40 N_VDD_c_40_p N_VSS_c_120_n 0.00106317f
cc_41 N_VDD_c_4_p N_VSS_c_121_n 0.00557569f
cc_42 N_VDD_c_4_p N_VSS_c_122_n 7.74609e-19
cc_43 N_VDD_c_7_p N_VSS_c_123_n 7.74609e-19
cc_44 N_VDD_c_16_p N_A_XI7.X0_CG 9.92565e-19
cc_45 N_VDD_XI7.X0_PGD N_A_c_171_n 3.90792e-19
cc_46 N_VDD_XI7.X0_PGD N_A_c_172_n 5.17967e-19
cc_47 N_VDD_c_4_p N_A_c_172_n 3.35498e-19
cc_48 N_VDD_c_7_p N_A_c_172_n 4.32724e-19
cc_49 N_VDD_c_15_p N_A_c_172_n 4.1682e-19
cc_50 N_VDD_c_16_p N_A_c_172_n 5.53168e-19
cc_51 N_VDD_c_11_p N_A_c_177_n 5.52801e-19
cc_52 N_VDD_c_12_p N_A_c_177_n 4.1541e-19
cc_53 N_VDD_c_31_p N_A_c_179_n 5.53687e-19
cc_54 N_VDD_c_31_p N_A_c_180_n 4.71537e-19
cc_55 N_VDD_XI6.X0_S N_BI_XI6.X0_D 3.43419e-19
cc_56 N_VDD_c_4_p N_BI_XI6.X0_D 3.70842e-19
cc_57 N_VDD_c_36_p N_BI_XI6.X0_D 3.72199e-19
cc_58 N_VDD_XI6.X0_S N_BI_c_253_n 3.48267e-19
cc_59 N_VDD_c_4_p N_BI_c_253_n 4.45573e-19
cc_60 N_VDD_c_36_p N_BI_c_253_n 5.2846e-19
cc_61 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_62 N_VDD_c_38_p N_AI_XI8.X0_D 3.72199e-19
cc_63 N_VDD_XI5.X0_PGD N_AI_XI2.X0_PGD 2.73831e-19
cc_64 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.86706e-19
cc_65 N_VDD_c_65_p N_AI_c_315_n 2.73831e-19
cc_66 N_VDD_c_66_p N_AI_c_316_n 2.86706e-19
cc_67 N_VDD_XI8.X0_S N_AI_c_317_n 3.48267e-19
cc_68 N_VDD_c_38_p N_AI_c_317_n 5.226e-19
cc_69 N_VDD_c_7_p N_AI_c_317_n 5.01863e-19
cc_70 N_VDD_c_15_p N_AI_c_320_n 0.00114922f
cc_71 N_VDD_c_7_p N_AI_c_321_n 2.39469e-19
cc_72 N_VDD_c_12_p N_B_XI5.X0_CG 0.00237871f
cc_73 N_VDD_XI5.X0_PGD N_B_c_359_n 3.9688e-19
cc_74 N_VDD_XI7.X0_PGD N_B_c_359_n 2.07132e-19
cc_75 N_VDD_c_31_p N_B_c_361_n 3.8625e-19
cc_76 N_VDD_c_11_p N_B_c_361_n 6.84022e-19
cc_77 N_VDD_c_12_p N_B_c_361_n 8.63725e-19
cc_78 N_VDD_c_11_p N_B_c_364_n 4.85469e-19
cc_79 N_VDD_c_12_p N_B_c_364_n 0.0014909f
cc_80 N_VDD_c_16_p N_B_c_364_n 5.33198e-19
cc_81 N_VSS_XI5.X0_D N_A_XI2.X0_S 3.43419e-19
cc_82 N_VSS_c_106_n N_A_c_182_n 0.00236445f
cc_83 N_VSS_XI8.X0_PGD N_A_c_171_n 3.86211e-19
cc_84 N_VSS_XI7.X0_S N_A_c_172_n 9.18655e-19
cc_85 N_VSS_c_97_n N_A_c_172_n 4.08476e-19
cc_86 N_VSS_c_98_n N_A_c_172_n 0.00149476f
cc_87 N_VSS_c_101_n N_A_c_172_n 2.91598e-19
cc_88 N_VSS_c_121_n N_A_c_172_n 2.51207e-19
cc_89 N_VSS_XI5.X0_D N_A_c_189_n 9.18655e-19
cc_90 N_VSS_c_97_n N_A_c_189_n 0.00202821f
cc_91 N_VSS_c_97_n N_A_c_177_n 0.0012307f
cc_92 N_VSS_c_135_p N_A_c_179_n 3.48564e-19
cc_93 N_VSS_c_93_n N_A_c_179_n 5.0102e-19
cc_94 N_VSS_c_106_n N_A_c_179_n 4.64764e-19
cc_95 N_VSS_c_110_n N_A_c_179_n 4.46304e-19
cc_96 N_VSS_c_93_n N_A_c_180_n 4.26083e-19
cc_97 N_VSS_c_102_n N_A_c_180_n 5.39888e-19
cc_98 N_VSS_c_106_n N_A_c_180_n 0.001324f
cc_99 N_VSS_XI5.X0_D N_BI_XI6.X0_D 3.43419e-19
cc_100 N_VSS_c_97_n N_BI_XI6.X0_D 3.48267e-19
cc_101 N_VSS_XI5.X0_D N_BI_c_253_n 3.48267e-19
cc_102 N_VSS_c_97_n N_BI_c_253_n 0.0010124f
cc_103 N_VSS_c_110_n N_BI_c_253_n 6.76595e-19
cc_104 N_VSS_c_121_n N_BI_c_253_n 6.07981e-19
cc_105 N_VSS_c_97_n N_BI_c_262_n 5.26238e-19
cc_106 N_VSS_c_121_n N_BI_c_262_n 7.0632e-19
cc_107 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_108 N_VSS_c_98_n N_AI_XI8.X0_D 3.48267e-19
cc_109 N_VSS_c_98_n N_AI_XI2.X0_PGD 2.04949e-19
cc_110 N_VSS_XI7.X0_S N_AI_c_317_n 3.48267e-19
cc_111 N_VSS_c_93_n N_AI_c_317_n 0.00173262f
cc_112 N_VSS_c_98_n N_AI_c_317_n 0.00129107f
cc_113 N_VSS_c_110_n N_AI_c_317_n 9.31051e-19
cc_114 N_VSS_c_98_n N_AI_c_320_n 0.00170897f
cc_115 N_VSS_c_98_n N_AI_c_330_n 2.82216e-19
cc_116 N_VSS_c_101_n N_AI_c_321_n 0.00934196f
cc_117 N_VSS_c_102_n N_B_XI6.X0_CG 9.70552e-19
cc_118 N_VSS_XI6.X0_PGD N_B_c_359_n 3.923e-19
cc_119 N_VSS_XI8.X0_PGD N_B_c_359_n 2.07132e-19
cc_120 N_VSS_c_110_n N_B_c_361_n 7.87668e-19
cc_121 N_VSS_c_97_n N_B_c_371_n 5.49592e-19
cc_122 N_VSS_c_101_n N_B_c_372_n 2.27662e-19
cc_123 N_VSS_XI7.X0_S N_C_XI4.X0_S 3.43419e-19
cc_124 N_VSS_c_98_n N_C_XI4.X0_S 3.48267e-19
cc_125 N_VSS_XI7.X0_S N_C_c_433_n 3.48267e-19
cc_126 N_VSS_c_98_n N_C_c_433_n 5.64614e-19
cc_127 N_A_c_199_p N_BI_XI2.X0_CG 2.16788e-19
cc_128 N_A_XI3.X0_PGD N_BI_c_265_n 8.79767e-19
cc_129 N_A_c_172_n N_BI_c_253_n 0.00115944f
cc_130 N_A_c_189_n N_BI_c_262_n 0.00163472f
cc_131 N_A_c_199_p N_BI_c_262_n 0.00112713f
cc_132 N_A_c_199_p N_BI_c_269_n 5.2034e-19
cc_133 N_A_c_189_n N_BI_c_270_n 3.37713e-19
cc_134 N_A_XI3.X0_PGD N_BI_c_271_n 0.00245019f
cc_135 N_A_c_207_p N_BI_c_271_n 3.56342e-19
cc_136 N_A_c_199_p N_BI_c_273_n 0.00124805f
cc_137 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174421f
cc_138 N_A_c_189_n N_AI_XI2.X0_PGD 8.48901e-19
cc_139 N_A_c_211_p N_AI_c_315_n 0.00195894f
cc_140 N_A_c_199_p N_AI_c_315_n 0.00178666f
cc_141 N_A_c_213_p N_AI_c_316_n 0.00202303f
cc_142 N_A_c_172_n N_AI_c_317_n 0.00165136f
cc_143 N_A_c_172_n N_AI_c_320_n 0.00201403f
cc_144 N_A_XI3.X0_PGD N_B_XI3.X0_CG 8.79767e-19
cc_145 N_A_c_207_p N_B_XI3.X0_CG 0.00234701f
cc_146 N_A_c_171_n N_B_c_359_n 0.0036024f
cc_147 N_A_c_172_n N_B_c_359_n 5.44634e-19
cc_148 N_A_c_180_n N_B_c_377_n 4.18059e-19
cc_149 N_A_c_172_n N_B_c_361_n 7.76373e-19
cc_150 N_A_c_189_n N_B_c_361_n 0.00128334f
cc_151 N_A_c_172_n N_B_c_380_n 3.26436e-19
cc_152 N_A_c_199_p N_B_c_381_n 3.96409e-19
cc_153 N_A_c_225_p N_B_c_381_n 9.9319e-19
cc_154 N_A_c_207_p N_B_c_381_n 4.87397e-19
cc_155 N_A_c_171_n N_B_c_364_n 3.81736e-19
cc_156 N_A_c_189_n N_B_c_364_n 5.63683e-19
cc_157 N_A_c_172_n N_B_c_386_n 3.8563e-19
cc_158 N_A_XI3.X0_PGD N_B_c_387_n 0.00312702f
cc_159 N_A_c_207_p N_B_c_387_n 0.00145837f
cc_160 N_A_c_189_n N_B_c_371_n 0.002414f
cc_161 N_A_c_233_p N_B_c_371_n 3.98537e-19
cc_162 N_A_c_199_p N_B_c_371_n 6.08993e-19
cc_163 N_A_c_172_n N_B_c_372_n 0.00197865f
cc_164 N_A_c_236_p N_C_c_435_n 2.22411e-19
cc_165 N_A_c_237_p N_C_c_436_n 4.03103e-19
cc_166 N_A_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_167 N_A_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_168 N_A_c_233_p N_Z_XI2.X0_D 3.48267e-19
cc_169 N_A_c_199_p N_Z_XI2.X0_D 9.18655e-19
cc_170 N_A_c_236_p N_Z_XI2.X0_D 3.48267e-19
cc_171 N_A_XI2.X0_S N_Z_c_463_n 3.48267e-19
cc_172 N_A_XI3.X0_S N_Z_c_463_n 3.48267e-19
cc_173 N_A_XI3.X0_PGD N_Z_c_463_n 5.57521e-19
cc_174 N_A_c_189_n N_Z_c_463_n 9.24e-19
cc_175 N_A_c_233_p N_Z_c_463_n 7.8992e-19
cc_176 N_A_c_199_p N_Z_c_463_n 0.00158543f
cc_177 N_A_c_236_p N_Z_c_463_n 8.08848e-19
cc_178 N_BI_XI2.X0_CG N_AI_XI2.X0_PGD 8.63152e-19
cc_179 N_BI_c_270_n N_AI_XI2.X0_PGD 0.00312702f
cc_180 N_BI_c_253_n N_AI_c_317_n 3.22835e-19
cc_181 N_BI_c_262_n N_AI_c_320_n 3.68388e-19
cc_182 N_BI_c_270_n N_AI_c_330_n 2.00604e-19
cc_183 N_BI_c_262_n N_B_c_361_n 0.00136623f
cc_184 N_BI_c_262_n N_B_c_380_n 6.77523e-19
cc_185 N_BI_c_270_n N_B_c_380_n 4.99367e-19
cc_186 N_BI_c_269_n N_B_c_381_n 0.00186236f
cc_187 N_BI_c_271_n N_B_c_381_n 4.99367e-19
cc_188 N_BI_c_273_n N_B_c_381_n 0.00166575f
cc_189 N_BI_c_270_n N_B_c_386_n 0.00513784f
cc_190 N_BI_c_271_n N_B_c_386_n 7.2092e-19
cc_191 N_BI_c_269_n N_B_c_387_n 4.99367e-19
cc_192 N_BI_c_270_n N_B_c_387_n 6.22265e-19
cc_193 N_BI_c_271_n N_B_c_387_n 0.00499463f
cc_194 N_BI_c_262_n N_B_c_371_n 0.00525284f
cc_195 N_BI_c_262_n N_B_c_405_n 2.67017e-19
cc_196 N_BI_c_273_n N_B_c_405_n 0.0013533f
cc_197 N_BI_c_293_p N_B_c_405_n 0.00340518f
cc_198 N_BI_c_262_n N_B_c_408_n 4.99817e-19
cc_199 N_BI_c_273_n N_B_c_408_n 9.35879e-19
cc_200 N_BI_c_296_p N_B_c_408_n 7.59935e-19
cc_201 N_BI_c_293_p N_B_c_411_n 0.00181541f
cc_202 N_BI_c_262_n N_B_c_412_n 0.00138818f
cc_203 N_BI_c_273_n N_B_c_412_n 8.23093e-19
cc_204 N_BI_c_262_n N_C_c_437_n 3.43796e-19
cc_205 N_BI_c_262_n N_C_c_436_n 7.49861e-19
cc_206 N_BI_c_269_n N_C_c_436_n 9.95458e-19
cc_207 N_BI_c_296_p N_C_c_436_n 3.37189e-19
cc_208 N_BI_c_262_n N_Z_c_463_n 0.00187303f
cc_209 N_BI_c_269_n N_Z_c_463_n 0.00192908f
cc_210 N_BI_c_270_n N_Z_c_463_n 8.66889e-19
cc_211 N_BI_c_271_n N_Z_c_463_n 8.66889e-19
cc_212 N_BI_c_273_n N_Z_c_463_n 7.39431e-19
cc_213 N_BI_c_293_p N_Z_c_463_n 0.00210701f
cc_214 N_BI_c_296_p N_Z_c_463_n 9.92397e-19
cc_215 N_AI_XI2.X0_PGD N_B_c_414_n 8.79767e-19
cc_216 N_AI_c_330_n N_B_c_414_n 0.00234701f
cc_217 N_AI_c_320_n N_B_c_380_n 5.22873e-19
cc_218 N_AI_c_330_n N_B_c_380_n 4.87397e-19
cc_219 N_AI_XI2.X0_PGD N_B_c_386_n 0.00312702f
cc_220 N_AI_c_320_n N_B_c_386_n 4.3265e-19
cc_221 N_AI_c_330_n N_B_c_386_n 0.00145837f
cc_222 N_AI_c_320_n N_B_c_372_n 0.00441104f
cc_223 N_AI_c_320_n N_B_c_405_n 3.85994e-19
cc_224 N_AI_c_320_n N_C_c_433_n 0.00187508f
cc_225 N_AI_c_317_n N_C_c_437_n 2.87718e-19
cc_226 N_AI_c_320_n N_C_c_437_n 8.98954e-19
cc_227 N_AI_c_320_n N_C_c_436_n 5.19511e-19
cc_228 N_AI_XI2.X0_PGD N_Z_c_463_n 2.98914e-19
cc_229 N_B_c_371_n N_C_c_433_n 8.83421e-19
cc_230 N_B_c_381_n N_C_c_436_n 9.42245e-19
cc_231 N_B_c_371_n N_C_c_436_n 2.24447e-19
cc_232 N_B_c_408_n N_C_c_436_n 0.00527131f
cc_233 N_B_c_380_n N_Z_c_463_n 0.00210511f
cc_234 N_B_c_381_n N_Z_c_463_n 0.00187303f
cc_235 N_B_c_387_n N_Z_c_463_n 8.66889e-19
cc_236 N_B_c_405_n N_Z_c_463_n 4.75654e-19
cc_237 N_C_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_238 N_C_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_239 N_C_c_433_n N_Z_XI4.X0_D 3.48267e-19
cc_240 N_C_c_435_n N_Z_XI4.X0_D 3.48267e-19
cc_241 N_C_XI4.X0_S N_Z_c_463_n 3.48267e-19
cc_242 N_C_XI1.X0_S N_Z_c_463_n 3.48267e-19
cc_243 N_C_c_433_n N_Z_c_463_n 5.74266e-19
cc_244 N_C_c_435_n N_Z_c_463_n 5.79289e-19
cc_245 N_C_c_436_n N_Z_c_463_n 4.30842e-19
*
.ends
*
*
.subckt MAJ3_HPNW4 A B C Y VDD VSS
xgate (VDD VSS A B C Y) G4_MAJ3_N1
.ends
*
* File: G3_MIN3_T6_N1.pex.netlist
* Created: Sun Apr 10 19:28:11 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MIN3_T6_N1_VSS 2 4 6 10 12 22 27 32 37 40 42 45 60 65 70 75 88 89
+ 93 99 102 103 108 Vss
c79 109 Vss 6.38121e-19
c80 108 Vss 0.00185802f
c81 103 Vss 0.00201533f
c82 99 Vss 0.0091126f
c83 94 Vss 0.00136513f
c84 93 Vss 0.00679427f
c85 89 Vss 6.52641e-19
c86 88 Vss 0.00390198f
c87 75 Vss 0.00302736f
c88 70 Vss 3.56438e-22
c89 65 Vss 0.00159414f
c90 60 Vss 9.05888e-19
c91 45 Vss 0.0850774f
c92 42 Vss 0.0849587f
c93 37 Vss 0.0679309f
c94 32 Vss 0.103393f
c95 27 Vss 0.306892f
c96 22 Vss 0.138043f
c97 12 Vss 0.00262003f
c98 10 Vss 0.0805405f
c99 6 Vss 0.0807339f
c100 4 Vss 0.00185192f
c101 2 Vss 0.0794633f
r102 107 108 3.66771
r103 103 107 0.655813
r104 100 109 0.494161
r105 100 102 12.1285
r106 99 108 0.652036
r107 99 102 0.87525
r108 95 109 0.128424
r109 93 109 0.494161
r110 93 94 10.0862
r111 88 94 0.652036
r112 87 89 0.655813
r113 87 88 9.08593
r114 70 103 1.82344
r115 65 95 4.33457
r116 60 75 1.16709
r117 60 89 1.82344
r118 45 47 1.8672
r119 42 44 1.8672
r120 40 75 0.50025
r121 37 40 1.92555
r122 33 47 0.0685365
r123 32 34 0.652036
r124 32 33 2.8008
r125 29 47 0.5835
r126 28 42 0.0685365
r127 27 45 0.0685365
r128 27 28 10.9698
r129 24 44 0.5835
r130 23 37 0.0685365
r131 22 44 0.0685365
r132 22 23 4.7847
r133 12 70 1.16709
r134 10 34 2.5674
r135 6 29 2.5674
r136 4 65 1.16709
r137 2 24 2.5674
.ends

.subckt PM_G3_MIN3_T6_N1_VDD 2 4 8 10 12 22 27 32 42 45 60 61 63 65 69 71 73 78
+ 81 83 Vss
c82 83 Vss 0.00427875f
c83 79 Vss 7.70868e-19
c84 78 Vss 0.00350656f
c85 73 Vss 0.00126506f
c86 71 Vss 0.0122742f
c87 69 Vss 0.00176475f
c88 65 Vss 0.00137661f
c89 63 Vss 7.01183e-19
c90 62 Vss 0.00177567f
c91 61 Vss 0.00769188f
c92 60 Vss 0.00512434f
c93 45 Vss 0.0848894f
c94 42 Vss 0.0854608f
c95 38 Vss 0.0711342f
c96 32 Vss 0.106688f
c97 27 Vss 0.309245f
c98 22 Vss 0.14138f
c99 12 Vss 0.0779484f
c100 10 Vss 0.0024321f
c101 8 Vss 0.0787627f
c102 4 Vss 0.0785563f
c103 2 Vss 0.00185192f
r104 78 81 0.349767
r105 77 78 3.66771
r106 73 81 0.306046
r107 73 75 1.82344
r108 72 79 0.494161
r109 71 77 0.652036
r110 71 72 13.0037
r111 67 79 0.128424
r112 67 69 4.33457
r113 65 83 1.16709
r114 63 65 1.82344
r115 61 79 0.494161
r116 61 62 10.0862
r117 60 63 0.655813
r118 59 62 0.652036
r119 59 60 9.08593
r120 45 46 1.8672
r121 42 43 1.8672
r122 38 83 0.50025
r123 38 40 1.92555
r124 33 45 0.0685365
r125 32 34 0.652036
r126 32 33 2.8008
r127 29 45 0.5835
r128 28 43 0.0685365
r129 27 46 0.0685365
r130 27 28 10.9698
r131 24 42 0.5835
r132 23 40 0.0685365
r133 22 42 0.0685365
r134 22 23 4.7847
r135 12 34 2.5674
r136 10 75 1.16709
r137 8 29 2.5674
r138 4 24 2.5674
r139 2 69 1.16709
.ends

.subckt PM_G3_MIN3_T6_N1_Z 2 4 6 8 48 56 59 61 Vss
c50 61 Vss 0.00482259f
c51 56 Vss 0.00183713f
c52 48 Vss 0.00151912f
c53 8 Vss 0.00176753f
c54 6 Vss 0.00171956f
c55 4 Vss 6.64706e-19
c56 2 Vss 6.16734e-19
r57 61 63 2.79246
r58 59 61 0.125036
r59 56 59 2.50071
r60 51 61 10.7364
r61 51 53 2.79246
r62 48 51 2.62575
r63 8 63 1.16709
r64 6 56 1.16709
r65 4 53 1.16709
r66 2 48 1.16709
.ends

.subckt PM_G3_MIN3_T6_N1_C 2 4 6 8 14 20 29 32 37 42 Vss
c31 42 Vss 0.0053281f
c32 37 Vss 0.00169525f
c33 32 Vss 0.00511278f
c34 29 Vss 5.02822e-19
c35 20 Vss 0.268178f
c36 14 Vss 0.269305f
r37 32 42 1.16709
r38 29 37 1.16709
r39 29 32 10.0654
r40 20 42 0.50025
r41 14 37 0.50025
r42 6 8 7.5855
r43 6 20 1.80885
r44 2 4 7.5855
r45 2 14 1.80885
.ends

.subckt PM_G3_MIN3_T6_N1_B 2 4 6 8 17 18 26 32 35 Vss
c28 35 Vss 0.00171406f
c29 32 Vss 3.1388e-19
c30 26 Vss 0.0844898f
c31 18 Vss 0.0345851f
c32 17 Vss 0.0963137f
c33 6 Vss 0.292132f
c34 2 Vss 0.340186f
r35 29 35 1.16709
r36 29 32 0.0729375
r37 24 35 0.0476429
r38 24 26 1.92555
r39 17 19 0.652036
r40 17 18 2.8008
r41 14 26 0.0685365
r42 13 18 0.652036
r43 6 8 7.5855
r44 6 19 2.5674
r45 4 14 2.5674
r46 2 4 7.5855
r47 2 13 2.5674
.ends

.subckt PM_G3_MIN3_T6_N1_A 2 4 6 8 29 34 37 41 46 Vss
c28 46 Vss 0.00547458f
c29 41 Vss 0.00144837f
c30 37 Vss 0.00108816f
c31 34 Vss 5.02933e-19
c32 29 Vss 3.18404e-19
c33 26 Vss 0.087104f
c34 6 Vss 0.296947f
c35 2 Vss 0.267858f
r36 37 46 1.16709
r37 34 37 0.0833571
r38 29 41 1.16709
r39 29 37 5.03269
r40 24 46 0.0476429
r41 24 26 1.92555
r42 19 26 0.0685365
r43 17 41 0.50025
r44 8 19 2.5674
r45 6 8 7.5855
r46 4 17 1.80885
r47 2 4 7.5855
.ends

.subckt G3_MIN3_T6_N1  VSS VDD Z C B A
*
* A	A
* B	B
* C	C
* Z	Z
* VDD	VDD
* VSS	VSS
XI9.X0 N_Z_XI9.X0_D N_VSS_XI9.X0_PGD N_C_XI9.X0_CG N_B_XI9.X0_PGS N_VDD_XI9.X0_S
+ TIGFET_HPNW4
XI6.X0 N_Z_XI6.X0_D N_VDD_XI6.X0_PGD N_C_XI6.X0_CG N_B_XI6.X0_PGS N_VSS_XI6.X0_S
+ TIGFET_HPNW4
XI11.X0 N_Z_XI11.X0_D N_VSS_XI11.X0_PGD N_A_XI11.X0_CG N_B_XI11.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW4
XI10.X0 N_Z_XI10.X0_D N_VDD_XI10.X0_PGD N_A_XI10.X0_CG N_B_XI10.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW4
XI8.X0 N_Z_XI11.X0_D N_VSS_XI8.X0_PGD N_C_XI8.X0_CG N_A_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI7.X0 N_Z_XI10.X0_D N_VDD_XI7.X0_PGD N_C_XI7.X0_CG N_A_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW4
*
x_PM_G3_MIN3_T6_N1_VSS N_VSS_XI9.X0_PGD N_VSS_XI6.X0_S N_VSS_XI11.X0_PGD
+ N_VSS_XI8.X0_PGD N_VSS_XI7.X0_S N_VSS_c_8_p N_VSS_c_24_p N_VSS_c_27_p
+ N_VSS_c_9_p N_VSS_c_15_p N_VSS_c_16_p N_VSS_c_61_p N_VSS_c_10_p N_VSS_c_2_p
+ N_VSS_c_6_p N_VSS_c_11_p N_VSS_c_12_p N_VSS_c_13_p N_VSS_c_19_p N_VSS_c_28_p
+ VSS N_VSS_c_31_p N_VSS_c_76_p Vss PM_G3_MIN3_T6_N1_VSS
x_PM_G3_MIN3_T6_N1_VDD N_VDD_XI9.X0_S N_VDD_XI6.X0_PGD N_VDD_XI10.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI7.X0_PGD N_VDD_c_87_n N_VDD_c_150_p N_VDD_c_160_p
+ N_VDD_c_153_p N_VDD_c_152_p N_VDD_c_88_n N_VDD_c_93_n N_VDD_c_99_n
+ N_VDD_c_100_n N_VDD_c_102_n N_VDD_c_105_n N_VDD_c_108_n N_VDD_c_142_p VDD
+ N_VDD_c_111_n Vss PM_G3_MIN3_T6_N1_VDD
x_PM_G3_MIN3_T6_N1_Z N_Z_XI9.X0_D N_Z_XI6.X0_D N_Z_XI11.X0_D N_Z_XI10.X0_D
+ N_Z_c_170_n N_Z_c_176_n Z N_Z_c_180_n Vss PM_G3_MIN3_T6_N1_Z
x_PM_G3_MIN3_T6_N1_C N_C_XI9.X0_CG N_C_XI6.X0_CG N_C_XI8.X0_CG N_C_XI7.X0_CG
+ N_C_c_212_n N_C_c_213_n C N_C_c_214_n N_C_c_215_n N_C_c_216_n Vss
+ PM_G3_MIN3_T6_N1_C
x_PM_G3_MIN3_T6_N1_B N_B_XI9.X0_PGS N_B_XI6.X0_PGS N_B_XI11.X0_PGS
+ N_B_XI10.X0_PGS N_B_c_247_n N_B_c_248_n N_B_c_256_n B N_B_c_258_n Vss
+ PM_G3_MIN3_T6_N1_B
x_PM_G3_MIN3_T6_N1_A N_A_XI11.X0_CG N_A_XI10.X0_CG N_A_XI8.X0_PGS N_A_XI7.X0_PGS
+ N_A_c_272_n A N_A_c_276_n N_A_c_282_n N_A_c_283_n Vss PM_G3_MIN3_T6_N1_A
cc_1 N_VSS_XI6.X0_S N_VDD_XI9.X0_S 4.21365e-19
cc_2 N_VSS_c_2_p N_VDD_XI9.X0_S 3.8999e-19
cc_3 N_VSS_XI9.X0_PGD N_VDD_XI6.X0_PGD 6.1888e-19
cc_4 N_VSS_XI11.X0_PGD N_VDD_XI10.X0_PGD 6.1888e-19
cc_5 N_VSS_XI7.X0_S N_VDD_XI8.X0_S 4.21365e-19
cc_6 N_VSS_c_6_p N_VDD_XI8.X0_S 3.8999e-19
cc_7 N_VSS_XI8.X0_PGD N_VDD_XI7.X0_PGD 5.98857e-19
cc_8 N_VSS_c_8_p N_VDD_c_87_n 6.35797e-19
cc_9 N_VSS_c_9_p N_VDD_c_88_n 2.61781e-19
cc_10 N_VSS_c_10_p N_VDD_c_88_n 0.00161042f
cc_11 N_VSS_c_11_p N_VDD_c_88_n 0.00118088f
cc_12 N_VSS_c_12_p N_VDD_c_88_n 0.00296683f
cc_13 N_VSS_c_13_p N_VDD_c_88_n 0.00183744f
cc_14 N_VSS_c_9_p N_VDD_c_93_n 9.27292e-19
cc_15 N_VSS_c_15_p N_VDD_c_93_n 3.72495e-19
cc_16 N_VSS_c_16_p N_VDD_c_93_n 8.87931e-19
cc_17 N_VSS_c_10_p N_VDD_c_93_n 9.0356e-19
cc_18 N_VSS_c_11_p N_VDD_c_93_n 4.3265e-19
cc_19 N_VSS_c_19_p N_VDD_c_93_n 3.0156e-19
cc_20 N_VSS_c_12_p N_VDD_c_99_n 0.00167687f
cc_21 N_VSS_c_10_p N_VDD_c_100_n 0.00121886f
cc_22 N_VSS_c_19_p N_VDD_c_100_n 3.71304e-19
cc_23 N_VSS_XI6.X0_S N_VDD_c_102_n 4.24828e-19
cc_24 N_VSS_c_24_p N_VDD_c_102_n 0.00115189f
cc_25 N_VSS_c_2_p N_VDD_c_102_n 4.59126e-19
cc_26 N_VSS_c_24_p N_VDD_c_105_n 9.72233e-19
cc_27 N_VSS_c_27_p N_VDD_c_105_n 8.14547e-19
cc_28 N_VSS_c_28_p N_VDD_c_105_n 3.32851e-19
cc_29 N_VSS_XI7.X0_S N_VDD_c_108_n 3.8999e-19
cc_30 N_VSS_c_6_p N_VDD_c_108_n 5.78716e-19
cc_31 N_VSS_c_31_p N_VDD_c_108_n 0.00180659f
cc_32 N_VSS_c_10_p N_VDD_c_111_n 3.8999e-19
cc_33 N_VSS_c_11_p N_VDD_c_111_n 0.00181085f
cc_34 N_VSS_c_10_p N_Z_XI9.X0_D 8.835e-19
cc_35 N_VSS_c_11_p N_Z_XI9.X0_D 0.00246958f
cc_36 N_VSS_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_37 N_VSS_c_2_p N_Z_XI6.X0_D 3.48267e-19
cc_38 N_VSS_XI6.X0_S N_Z_XI10.X0_D 3.43419e-19
cc_39 N_VSS_XI7.X0_S N_Z_XI10.X0_D 3.43419e-19
cc_40 N_VSS_c_2_p N_Z_XI10.X0_D 3.48267e-19
cc_41 N_VSS_c_6_p N_Z_XI10.X0_D 3.48267e-19
cc_42 N_VSS_XI6.X0_S N_Z_c_170_n 3.48267e-19
cc_43 N_VSS_c_10_p N_Z_c_170_n 0.00217565f
cc_44 N_VSS_c_2_p N_Z_c_170_n 5.69026e-19
cc_45 N_VSS_c_11_p N_Z_c_170_n 8.835e-19
cc_46 N_VSS_c_12_p N_Z_c_170_n 7.10715e-19
cc_47 N_VSS_c_19_p N_Z_c_170_n 3.30259e-19
cc_48 N_VSS_XI6.X0_S N_Z_c_176_n 3.48267e-19
cc_49 N_VSS_XI7.X0_S N_Z_c_176_n 3.48267e-19
cc_50 N_VSS_c_2_p N_Z_c_176_n 5.69026e-19
cc_51 N_VSS_c_6_p N_Z_c_176_n 5.69026e-19
cc_52 N_VSS_c_2_p N_Z_c_180_n 0.00191849f
cc_53 N_VSS_c_12_p N_Z_c_180_n 5.57576e-19
cc_54 N_VSS_c_19_p N_Z_c_180_n 0.00201399f
cc_55 N_VSS_c_28_p N_Z_c_180_n 5.26184e-19
cc_56 N_VSS_XI9.X0_PGD N_C_c_212_n 4.30517e-19
cc_57 N_VSS_XI8.X0_PGD N_C_c_213_n 5.02359e-19
cc_58 N_VSS_c_28_p N_C_c_214_n 2.73385e-19
cc_59 N_VSS_XI9.X0_PGD N_C_c_215_n 4.3583e-19
cc_60 N_VSS_XI8.X0_PGD N_C_c_216_n 3.76133e-19
cc_61 N_VSS_c_61_p N_C_c_216_n 2.17009e-19
cc_62 N_VSS_XI9.X0_PGD N_B_XI9.X0_PGS 0.00109504f
cc_63 N_VSS_XI11.X0_PGD N_B_XI9.X0_PGS 2.15671e-19
cc_64 N_VSS_XI11.X0_PGD N_B_XI11.X0_PGS 0.00177732f
cc_65 N_VSS_XI8.X0_PGD N_B_XI11.X0_PGS 2.22194e-19
cc_66 N_VSS_c_61_p N_B_c_247_n 0.00177732f
cc_67 N_VSS_c_24_p N_B_c_248_n 0.00731987f
cc_68 N_VSS_c_16_p N_B_c_248_n 0.00109504f
cc_69 N_VSS_c_2_p B 2.11465e-19
cc_70 N_VSS_c_12_p B 2.74582e-19
cc_71 N_VSS_c_19_p B 2.99651e-19
cc_72 N_VSS_c_24_p N_A_XI11.X0_CG 2.66861e-19
cc_73 N_VSS_c_2_p N_A_c_272_n 3.13396e-19
cc_74 N_VSS_c_28_p N_A_c_272_n 5.88825e-19
cc_75 N_VSS_c_28_p A 5.88825e-19
cc_76 N_VSS_c_76_p A 2.39495e-19
cc_77 N_VSS_c_2_p N_A_c_276_n 0.00159849f
cc_78 N_VSS_c_28_p N_A_c_276_n 0.00924443f
cc_79 N_VSS_c_76_p N_A_c_276_n 5.12768e-19
cc_80 N_VDD_XI9.X0_S N_Z_XI9.X0_D 3.43419e-19
cc_81 N_VDD_c_93_n N_Z_XI9.X0_D 4.3265e-19
cc_82 N_VDD_c_102_n N_Z_XI9.X0_D 3.48267e-19
cc_83 N_VDD_c_100_n N_Z_XI6.X0_D 9.44213e-19
cc_84 N_VDD_c_111_n N_Z_XI6.X0_D 0.00246958f
cc_85 N_VDD_XI9.X0_S N_Z_XI11.X0_D 3.43419e-19
cc_86 N_VDD_XI8.X0_S N_Z_XI11.X0_D 3.43419e-19
cc_87 N_VDD_c_102_n N_Z_XI11.X0_D 3.48267e-19
cc_88 N_VDD_c_105_n N_Z_XI11.X0_D 4.3265e-19
cc_89 N_VDD_c_108_n N_Z_XI11.X0_D 3.72199e-19
cc_90 N_VDD_XI9.X0_S N_Z_c_170_n 3.48267e-19
cc_91 N_VDD_c_88_n N_Z_c_170_n 0.0013145f
cc_92 N_VDD_c_93_n N_Z_c_170_n 7.37531e-19
cc_93 N_VDD_c_100_n N_Z_c_170_n 0.00186578f
cc_94 N_VDD_c_102_n N_Z_c_170_n 7.73813e-19
cc_95 N_VDD_c_111_n N_Z_c_170_n 8.835e-19
cc_96 N_VDD_XI9.X0_S N_Z_c_176_n 3.48267e-19
cc_97 N_VDD_XI8.X0_S N_Z_c_176_n 3.48267e-19
cc_98 N_VDD_c_102_n N_Z_c_176_n 8.00908e-19
cc_99 N_VDD_c_105_n N_Z_c_176_n 5.78499e-19
cc_100 N_VDD_c_108_n N_Z_c_176_n 8.53368e-19
cc_101 N_VDD_c_93_n N_Z_c_180_n 8.36802e-19
cc_102 N_VDD_c_88_n C 2.63478e-19
cc_103 N_VDD_c_93_n C 0.00145322f
cc_104 N_VDD_c_102_n C 0.00155931f
cc_105 N_VDD_c_88_n N_C_c_214_n 2.14517e-19
cc_106 N_VDD_c_93_n N_C_c_214_n 8.61717e-19
cc_107 N_VDD_c_102_n N_C_c_214_n 0.00183615f
cc_108 N_VDD_c_105_n N_C_c_214_n 0.00557625f
cc_109 N_VDD_c_142_p N_C_c_214_n 5.42852e-19
cc_110 N_VDD_c_93_n N_C_c_215_n 7.51813e-19
cc_111 N_VDD_c_102_n N_C_c_215_n 8.66889e-19
cc_112 N_VDD_c_102_n N_C_c_216_n 2.22969e-19
cc_113 N_VDD_c_105_n N_C_c_216_n 2.63125e-19
cc_114 N_VDD_c_142_p N_C_c_216_n 3.66936e-19
cc_115 N_VDD_XI6.X0_PGD N_B_XI9.X0_PGS 0.00135245f
cc_116 N_VDD_XI10.X0_PGD N_B_XI9.X0_PGS 4.12959e-19
cc_117 N_VDD_c_150_p N_B_XI11.X0_PGS 0.00109105f
cc_118 N_VDD_c_150_p N_B_c_256_n 0.00258419f
cc_119 N_VDD_c_152_p N_B_c_256_n 4.12959e-19
cc_120 N_VDD_c_153_p N_B_c_258_n 0.00495207f
cc_121 N_VDD_c_111_n N_B_c_258_n 4.60491e-19
cc_122 N_VDD_XI10.X0_PGD N_A_XI11.X0_CG 4.83278e-19
cc_123 N_VDD_XI7.X0_PGD N_A_XI8.X0_PGS 0.00141985f
cc_124 N_VDD_c_105_n N_A_XI8.X0_PGS 2.26738e-19
cc_125 N_VDD_XI10.X0_PGD N_A_c_282_n 5.50272e-19
cc_126 N_VDD_XI7.X0_PGD N_A_c_283_n 3.23173e-19
cc_127 N_VDD_c_160_p N_A_c_283_n 0.00145458f
cc_128 N_VDD_c_152_p N_A_c_283_n 2.17009e-19
cc_129 N_Z_c_170_n N_C_c_212_n 6.18749e-19
cc_130 N_Z_c_176_n N_C_c_213_n 8.38264e-19
cc_131 N_Z_c_180_n N_C_c_214_n 0.0071108f
cc_132 N_Z_c_176_n N_A_XI11.X0_CG 2.49716e-19
cc_133 N_Z_c_176_n N_A_c_276_n 3.55289e-19
cc_134 N_Z_c_180_n N_A_c_276_n 0.00276659f
cc_135 N_C_c_212_n N_B_XI9.X0_PGS 0.00830899f
cc_136 N_C_c_215_n N_B_XI9.X0_PGS 3.76133e-19
cc_137 N_C_c_212_n N_B_XI11.X0_PGS 8.90713e-19
cc_138 N_C_c_213_n N_B_XI11.X0_PGS 5.42381e-19
cc_139 N_C_c_215_n N_B_c_258_n 3.15193e-19
cc_140 N_C_c_213_n N_A_XI11.X0_CG 0.0020589f
cc_141 N_C_c_213_n N_A_XI8.X0_PGS 0.00810452f
cc_142 N_C_c_214_n N_A_c_276_n 0.00121525f
cc_143 N_C_c_216_n N_A_c_283_n 3.16599e-19
cc_144 N_B_XI9.X0_PGS N_A_XI11.X0_CG 0.00106357f
cc_145 N_B_XI11.X0_PGS N_A_XI11.X0_CG 0.00765248f
cc_146 B N_A_c_272_n 3.39698e-19
cc_147 N_B_c_258_n N_A_c_272_n 3.48267e-19
cc_148 B N_A_c_282_n 3.48267e-19
cc_149 N_B_c_258_n N_A_c_282_n 5.15124e-19
*
.ends
*
*
.subckt MIN3_HPNW4 A B C Y VDD VSS
xgate (VSS VDD Y C B A) G3_MIN3_T6_N1
.ends
*
* File: G4_MUX2_N1.pex.netlist
* Created: Wed Mar  9 17:10:36 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MUX2_N1_VDD 2 4 6 8 10 12 14 18 20 38 49 58 84 85 87 89 93 95 96
+ 99 101 105 107 111 113 115 120 122 124 125 126 127 128 134 139 148 Vss
c140 148 Vss 0.00577129f
c141 139 Vss 0.00441689f
c142 134 Vss 0.00586273f
c143 128 Vss 3.56526e-19
c144 127 Vss 2.39889e-19
c145 126 Vss 4.22747e-19
c146 125 Vss 2.39889e-19
c147 122 Vss 0.00188211f
c148 120 Vss 0.00629792f
c149 115 Vss 0.00178287f
c150 113 Vss 0.00614865f
c151 111 Vss 6.94069e-19
c152 107 Vss 0.00775764f
c153 105 Vss 0.001258f
c154 101 Vss 0.00169538f
c155 99 Vss 4.33371e-19
c156 96 Vss 6.1175e-19
c157 95 Vss 0.00337348f
c158 93 Vss 0.00135966f
c159 89 Vss 0.00148319f
c160 87 Vss 0.00118366f
c161 85 Vss 0.00653402f
c162 84 Vss 0.00317212f
c163 83 Vss 0.00175227f
c164 59 Vss 0.0798032f
c165 58 Vss 0.102888f
c166 49 Vss 0.0346129f
c167 48 Vss 0.100303f
c168 39 Vss 0.0355046f
c169 38 Vss 0.100457f
c170 20 Vss 0.00271849f
c171 18 Vss 0.0807095f
c172 14 Vss 0.0816769f
c173 12 Vss 0.00155055f
c174 10 Vss 0.0815741f
c175 8 Vss 0.0807057f
c176 6 Vss 0.0842982f
c177 4 Vss 0.0825471f
c178 2 Vss 0.00231862f
r179 121 128 0.551426
r180 121 122 4.16786
r181 120 128 0.551426
r182 119 120 13.3371
r183 115 128 0.0828784
r184 115 117 1.82344
r185 114 127 0.494161
r186 113 119 0.652036
r187 113 114 10.1279
r188 111 148 1.16709
r189 109 127 0.128424
r190 109 111 2.16729
r191 108 126 0.494161
r192 107 122 0.652036
r193 107 108 13.0037
r194 103 126 0.128424
r195 103 105 4.83471
r196 102 125 0.494161
r197 101 127 0.494161
r198 101 102 4.58464
r199 99 139 1.16709
r200 97 125 0.128424
r201 97 99 2.16729
r202 95 126 0.494161
r203 95 96 7.46046
r204 93 134 1.16709
r205 91 96 0.652036
r206 91 93 2.16729
r207 87 89 1.82344
r208 86 124 0.326018
r209 85 125 0.494161
r210 85 86 10.1279
r211 84 87 0.655813
r212 83 124 0.326018
r213 83 84 4.16786
r214 64 148 0.238214
r215 64 66 1.92555
r216 59 66 0.5835
r217 58 60 0.652036
r218 58 59 2.8008
r219 55 66 0.0685365
r220 51 139 0.238214
r221 49 51 1.45875
r222 48 52 0.652036
r223 48 51 1.45875
r224 45 49 0.652036
r225 41 134 0.238214
r226 39 41 1.45875
r227 38 42 0.652036
r228 38 41 1.45875
r229 35 39 0.652036
r230 20 117 1.16709
r231 18 60 2.5674
r232 14 55 2.5674
r233 12 105 1.16709
r234 10 52 2.5674
r235 8 45 2.5674
r236 6 35 2.5674
r237 4 42 2.5674
r238 2 89 1.16709
.ends

.subckt PM_G4_MUX2_N1_VSS 2 4 6 8 10 12 16 18 20 38 39 48 49 51 59 84 89 94 99
+ 104 109 118 123 132 141 142 146 152 153 158 164 170 172 177 179 181 182 183
+ 184 185 Vss
c132 185 Vss 4.28045e-19
c133 184 Vss 3.62111e-19
c134 183 Vss 3.87529e-19
c135 182 Vss 3.75522e-19
c136 179 Vss 0.00396469f
c137 177 Vss 0.00140343f
c138 172 Vss 0.00128299f
c139 170 Vss 0.00250671f
c140 164 Vss 0.00572414f
c141 158 Vss 0.00417852f
c142 153 Vss 5.94991e-19
c143 152 Vss 0.00253786f
c144 146 Vss 0.00510722f
c145 142 Vss 0.00100335f
c146 141 Vss 0.00361314f
c147 132 Vss 0.00636077f
c148 123 Vss 0.00367258f
c149 118 Vss 0.0040616f
c150 109 Vss 3.31973e-19
c151 104 Vss 0.00116949f
c152 99 Vss 0.00135225f
c153 94 Vss 3.56537e-19
c154 89 Vss 8.02281e-19
c155 84 Vss 0.00135359f
c156 65 Vss 0.0785271f
c157 59 Vss 0.0340359f
c158 58 Vss 0.0688517f
c159 49 Vss 0.0338093f
c160 48 Vss 0.0993447f
c161 39 Vss 0.0341976f
c162 38 Vss 0.0984533f
c163 20 Vss 0.0819076f
c164 18 Vss 0.00227065f
c165 16 Vss 0.0807095f
c166 12 Vss 0.0827078f
c167 10 Vss 0.0826808f
c168 8 Vss 0.00150258f
c169 6 Vss 0.00290641f
c170 4 Vss 0.081612f
c171 2 Vss 0.0842992f
r172 178 185 0.551426
r173 178 179 13.3371
r174 177 185 0.551426
r175 176 177 4.16786
r176 172 185 0.0828784
r177 171 184 0.494161
r178 170 179 0.652036
r179 170 171 4.41793
r180 166 184 0.128424
r181 165 183 0.494161
r182 164 176 0.652036
r183 164 165 13.0037
r184 160 183 0.128424
r185 159 182 0.494161
r186 158 184 0.494161
r187 158 159 10.2946
r188 154 182 0.128424
r189 152 183 0.494161
r190 152 153 7.46046
r191 148 153 0.652036
r192 147 181 0.326018
r193 146 182 0.494161
r194 146 147 10.1279
r195 141 181 0.326018
r196 140 142 0.655813
r197 140 141 4.16786
r198 109 172 1.82344
r199 104 132 1.16709
r200 104 166 2.16729
r201 99 160 4.83471
r202 94 123 1.16709
r203 94 154 2.16729
r204 89 118 1.16709
r205 89 148 2.16729
r206 84 142 1.82344
r207 65 132 0.238214
r208 63 65 1.8672
r209 60 63 0.0685365
r210 58 63 0.5835
r211 58 59 2.8008
r212 55 59 0.652036
r213 51 123 0.238214
r214 49 51 1.45875
r215 48 52 0.652036
r216 48 51 1.45875
r217 45 49 0.652036
r218 41 118 0.238214
r219 39 41 1.45875
r220 38 42 0.652036
r221 38 41 1.45875
r222 35 39 0.652036
r223 20 60 2.5674
r224 18 109 1.16709
r225 16 55 2.5674
r226 12 52 2.5674
r227 10 45 2.5674
r228 8 99 1.16709
r229 6 84 1.16709
r230 4 42 2.5674
r231 2 35 2.5674
.ends

.subckt PM_G4_MUX2_N1_ZI 2 4 6 8 28 50 55 60 65 81 82 91 Vss
c67 82 Vss 9.74571e-19
c68 81 Vss 0.00289684f
c69 65 Vss 0.00556163f
c70 60 Vss 8.37584e-19
c71 55 Vss 0.00123466f
c72 50 Vss 0.00178991f
c73 28 Vss 0.206432f
c74 23 Vss 0.0247918f
c75 8 Vss 0.00143442f
c76 6 Vss 0.00143442f
c77 4 Vss 0.0815973f
c78 2 Vss 0.0715834f
r79 87 91 0.494161
r80 83 91 0.494161
r81 81 91 0.128424
r82 81 82 13.2121
r83 77 82 0.652036
r84 60 87 3.66771
r85 55 83 4.33457
r86 50 65 1.16709
r87 50 77 2.16729
r88 31 65 0.0476429
r89 29 31 0.326018
r90 29 31 0.1167
r91 28 32 0.652036
r92 28 31 6.7686
r93 27 65 0.357321
r94 23 31 0.326018
r95 23 27 0.40845
r96 8 60 1.16709
r97 6 55 1.16709
r98 4 32 2.5674
r99 2 27 2.15895
.ends

.subckt PM_G4_MUX2_N1_Z 2 18 Vss
c12 18 Vss 2.88294e-19
c13 2 Vss 0.00150258f
r14 2 18 1.16709
.ends

.subckt PM_G4_MUX2_N1_SELI 2 6 8 21 33 35 36 38 43 53 58 72 77 78 Vss
c81 78 Vss 6.39942e-19
c82 77 Vss 5.11483e-19
c83 72 Vss 0.00145166f
c84 58 Vss 0.0021541f
c85 53 Vss 0.00198421f
c86 43 Vss 9.80359e-19
c87 38 Vss 0.00153196f
c88 36 Vss 2.15854e-19
c89 35 Vss 0.00258645f
c90 33 Vss 0.00238155f
c91 21 Vss 0.0575125f
c92 6 Vss 0.0575499f
c93 2 Vss 0.00172036f
r94 77 78 0.655813
r95 76 77 3.501
r96 72 76 0.655813
r97 43 53 1.16709
r98 43 72 2.00578
r99 43 46 0.833571
r100 38 58 1.16709
r101 38 78 2.00578
r102 35 46 0.0685365
r103 35 36 7.46046
r104 31 36 0.652036
r105 31 33 5.58493
r106 21 58 0.50025
r107 18 53 0.50025
r108 8 21 1.80885
r109 6 18 1.80885
r110 2 33 1.16709
.ends

.subckt PM_G4_MUX2_N1_SEL 2 4 6 8 16 17 22 26 37 40 41 44 45 46 47 52 58 63 68
+ 73 Vss
c78 73 Vss 0.00176698f
c79 68 Vss 0.00182856f
c80 63 Vss 0.00250521f
c81 58 Vss 7.07944e-19
c82 52 Vss 2.9409e-19
c83 47 Vss 2.03369e-19
c84 46 Vss 3.54223e-19
c85 45 Vss 7.77909e-19
c86 44 Vss 0.00151239f
c87 41 Vss 0.00163463f
c88 37 Vss 0.00192905f
c89 26 Vss 0.0575125f
c90 22 Vss 0.0712295f
c91 20 Vss 0.0247918f
c92 17 Vss 0.0358042f
c93 16 Vss 0.175331f
c94 8 Vss 0.0575125f
c95 2 Vss 0.084915f
r96 58 73 1.16709
r97 58 60 0.5835
r98 55 68 1.16709
r99 52 55 0.5835
r100 50 63 1.16709
r101 47 50 0.5835
r102 45 60 0.0685365
r103 45 46 1.70882
r104 43 46 0.652036
r105 43 44 2.50071
r106 42 52 0.0685365
r107 41 44 0.652036
r108 41 42 1.70882
r109 38 47 0.0685365
r110 38 40 1.62546
r111 37 52 0.0685365
r112 37 40 2.95918
r113 36 63 0.0476429
r114 33 73 0.50025
r115 26 68 0.50025
r116 22 63 0.357321
r117 20 36 0.326018
r118 20 22 0.40845
r119 17 36 6.7686
r120 16 36 0.326018
r121 16 36 0.1167
r122 13 17 0.652036
r123 8 33 1.80885
r124 6 26 1.80885
r125 4 22 2.15895
r126 2 13 2.5674
.ends

.subckt PM_G4_MUX2_N1_B 2 4 14 20 23 Vss
c31 23 Vss 0.00482401f
c32 20 Vss 4.63929e-19
c33 14 Vss 0.0843809f
c34 2 Vss 0.446304f
r35 17 23 1.16709
r36 17 20 0.0364688
r37 14 23 0.238214
r38 11 14 1.92555
r39 7 11 0.0685365
r40 4 7 2.5674
r41 2 4 12.837
.ends

.subckt PM_G4_MUX2_N1_A 2 4 14 20 23 Vss
c25 23 Vss 0.00557714f
c26 20 Vss 2.81445e-19
c27 14 Vss 0.0830192f
c28 2 Vss 0.44929f
r29 17 23 1.16709
r30 17 20 0.0729375
r31 12 23 0.238214
r32 12 14 1.92555
r33 7 14 0.0685365
r34 2 4 12.837
r35 2 7 2.5674
.ends

.subckt G4_MUX2_N1  VDD VSS Z SEL B A
*
* A	A
* B	B
* SEL	SEL
* Z	Z
* VSS	VSS
* VDD	VDD
XI7.X0 N_VDD_XI7.X0_D N_VSS_XI7.X0_PGD N_ZI_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_Z_XI7.X0_S TIGFET_HPNW4
XI1.X0 N_SELI_XI1.X0_D N_VDD_XI1.X0_PGD N_SEL_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI6.X0 N_Z_XI7.X0_S N_VDD_XI6.X0_PGD N_ZI_XI6.X0_CG N_VDD_XI6.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW4
XI2.X0 N_SELI_XI1.X0_D N_VSS_XI2.X0_PGD N_SEL_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI5.X0 N_ZI_XI5.X0_D N_VDD_XI5.X0_PGD N_SELI_XI5.X0_CG N_B_XI5.X0_PGS
+ N_VSS_XI6.X0_S TIGFET_HPNW4
XI3.X0 N_ZI_XI3.X0_D N_VSS_XI3.X0_PGD N_SEL_XI3.X0_CG N_B_XI3.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI4.X0 N_ZI_XI5.X0_D N_VDD_XI4.X0_PGD N_SEL_XI4.X0_CG N_A_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW4
XI0.X0 N_ZI_XI3.X0_D N_VSS_XI0.X0_PGD N_SELI_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW4
*
x_PM_G4_MUX2_N1_VDD N_VDD_XI7.X0_D N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS
+ N_VDD_XI6.X0_PGD N_VDD_XI6.X0_PGS N_VDD_XI2.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_14_p N_VDD_c_11_p N_VDD_c_136_p
+ N_VDD_c_18_p N_VDD_c_12_p N_VDD_c_46_p N_VDD_c_17_p N_VDD_c_22_p N_VDD_c_15_p
+ N_VDD_c_48_p N_VDD_c_20_p N_VDD_c_3_p N_VDD_c_6_p N_VDD_c_16_p N_VDD_c_28_p
+ N_VDD_c_8_p N_VDD_c_34_p N_VDD_c_9_p N_VDD_c_32_p VDD N_VDD_c_51_p
+ N_VDD_c_55_p N_VDD_c_58_p N_VDD_c_65_p N_VDD_c_25_p N_VDD_c_21_p N_VDD_c_95_p
+ Vss PM_G4_MUX2_N1_VDD
x_PM_G4_MUX2_N1_VSS N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS N_VSS_XI1.X0_S
+ N_VSS_XI6.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS N_VSS_XI3.X0_PGD
+ N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_151_n N_VSS_c_153_n N_VSS_c_265_p
+ N_VSS_c_154_n N_VSS_c_257_p N_VSS_c_156_n N_VSS_c_157_n N_VSS_c_158_n
+ N_VSS_c_162_n N_VSS_c_166_n N_VSS_c_170_n N_VSS_c_173_n N_VSS_c_176_n
+ N_VSS_c_180_n N_VSS_c_184_n N_VSS_c_185_n N_VSS_c_186_n N_VSS_c_187_n
+ N_VSS_c_189_n N_VSS_c_192_n N_VSS_c_193_n N_VSS_c_196_n N_VSS_c_199_n
+ N_VSS_c_200_n N_VSS_c_201_n N_VSS_c_202_n VSS N_VSS_c_206_n N_VSS_c_207_n
+ N_VSS_c_208_n N_VSS_c_209_n Vss PM_G4_MUX2_N1_VSS
x_PM_G4_MUX2_N1_ZI N_ZI_XI7.X0_CG N_ZI_XI6.X0_CG N_ZI_XI5.X0_D N_ZI_XI3.X0_D
+ N_ZI_c_278_n N_ZI_c_294_n N_ZI_c_280_n N_ZI_c_282_n N_ZI_c_287_n N_ZI_c_288_n
+ N_ZI_c_311_n N_ZI_c_326_p Vss PM_G4_MUX2_N1_ZI
x_PM_G4_MUX2_N1_Z N_Z_XI7.X0_S Z Vss PM_G4_MUX2_N1_Z
x_PM_G4_MUX2_N1_SELI N_SELI_XI1.X0_D N_SELI_XI5.X0_CG N_SELI_XI0.X0_CG
+ N_SELI_c_371_n N_SELI_c_356_n N_SELI_c_359_n N_SELI_c_387_n N_SELI_c_364_n
+ N_SELI_c_365_n N_SELI_c_367_n N_SELI_c_379_n N_SELI_c_381_n N_SELI_c_395_n
+ N_SELI_c_398_n Vss PM_G4_MUX2_N1_SELI
x_PM_G4_MUX2_N1_SEL N_SEL_XI1.X0_CG N_SEL_XI2.X0_CG N_SEL_XI3.X0_CG
+ N_SEL_XI4.X0_CG N_SEL_c_434_n N_SEL_c_460_n N_SEL_c_449_n N_SEL_c_495_p
+ N_SEL_c_436_n SEL N_SEL_c_438_n N_SEL_c_439_n N_SEL_c_440_n N_SEL_c_465_n
+ N_SEL_c_453_n N_SEL_c_468_n N_SEL_c_442_n N_SEL_c_443_n N_SEL_c_444_n
+ N_SEL_c_445_n Vss PM_G4_MUX2_N1_SEL
x_PM_G4_MUX2_N1_B N_B_XI5.X0_PGS N_B_XI3.X0_PGS N_B_c_518_n B N_B_c_514_n Vss
+ PM_G4_MUX2_N1_B
x_PM_G4_MUX2_N1_A N_A_XI4.X0_PGS N_A_XI0.X0_PGS N_A_c_544_n A N_A_c_550_n Vss
+ PM_G4_MUX2_N1_A
cc_1 N_VDD_XI1.X0_PGS N_VSS_XI7.X0_PGD 2.27468e-19
cc_2 N_VDD_XI6.X0_PGD N_VSS_XI7.X0_PGS 0.00173038f
cc_3 N_VDD_c_3_p N_VSS_XI6.X0_S 3.7884e-19
cc_4 N_VDD_XI1.X0_PGD N_VSS_XI2.X0_PGD 0.0016786f
cc_5 N_VDD_XI6.X0_PGS N_VSS_XI2.X0_PGS 2.11937e-19
cc_6 N_VDD_c_6_p N_VSS_XI2.X0_PGS 2.56778e-19
cc_7 N_VDD_XI5.X0_PGD N_VSS_XI3.X0_PGD 2.1536e-19
cc_8 N_VDD_c_8_p N_VSS_XI4.X0_S 3.7884e-19
cc_9 N_VDD_c_9_p N_VSS_XI4.X0_S 9.5668e-19
cc_10 N_VDD_XI4.X0_PGD N_VSS_XI0.X0_PGD 2.1536e-19
cc_11 N_VDD_c_11_p N_VSS_c_151_n 0.00173038f
cc_12 N_VDD_c_12_p N_VSS_c_151_n 3.60588e-19
cc_13 N_VDD_c_12_p N_VSS_c_153_n 3.80388e-19
cc_14 N_VDD_c_14_p N_VSS_c_154_n 0.0016786f
cc_15 N_VDD_c_15_p N_VSS_c_154_n 2.72324e-19
cc_16 N_VDD_c_16_p N_VSS_c_156_n 8.01165e-19
cc_17 N_VDD_c_17_p N_VSS_c_157_n 9.30123e-19
cc_18 N_VDD_c_18_p N_VSS_c_158_n 8.69498e-19
cc_19 N_VDD_c_12_p N_VSS_c_158_n 0.00141228f
cc_20 N_VDD_c_20_p N_VSS_c_158_n 8.51944e-19
cc_21 N_VDD_c_21_p N_VSS_c_158_n 3.48267e-19
cc_22 N_VDD_c_22_p N_VSS_c_162_n 8.56577e-19
cc_23 N_VDD_c_15_p N_VSS_c_162_n 0.00141228f
cc_24 N_VDD_c_6_p N_VSS_c_162_n 0.00181129f
cc_25 N_VDD_c_25_p N_VSS_c_162_n 3.48267e-19
cc_26 N_VDD_c_20_p N_VSS_c_166_n 3.92901e-19
cc_27 N_VDD_c_3_p N_VSS_c_166_n 4.58491e-19
cc_28 N_VDD_c_28_p N_VSS_c_166_n 7.06793e-19
cc_29 N_VDD_c_9_p N_VSS_c_166_n 2.71563e-19
cc_30 N_VDD_c_6_p N_VSS_c_170_n 2.93442e-19
cc_31 N_VDD_c_16_p N_VSS_c_170_n 0.00161703f
cc_32 N_VDD_c_32_p N_VSS_c_170_n 4.6996e-19
cc_33 N_VDD_c_8_p N_VSS_c_173_n 4.73473e-19
cc_34 N_VDD_c_34_p N_VSS_c_173_n 2.13058e-19
cc_35 N_VDD_c_9_p N_VSS_c_173_n 0.00165395f
cc_36 N_VDD_c_18_p N_VSS_c_176_n 3.66936e-19
cc_37 N_VDD_c_12_p N_VSS_c_176_n 0.00112249f
cc_38 N_VDD_c_20_p N_VSS_c_176_n 3.99794e-19
cc_39 N_VDD_c_21_p N_VSS_c_176_n 8.07896e-19
cc_40 N_VDD_c_22_p N_VSS_c_180_n 3.82294e-19
cc_41 N_VDD_c_15_p N_VSS_c_180_n 0.00112249f
cc_42 N_VDD_c_6_p N_VSS_c_180_n 9.55349e-19
cc_43 N_VDD_c_25_p N_VSS_c_180_n 8.0279e-19
cc_44 N_VDD_c_16_p N_VSS_c_184_n 2.03837e-19
cc_45 N_VDD_c_22_p N_VSS_c_185_n 3.85245e-19
cc_46 N_VDD_c_46_p N_VSS_c_186_n 4.93614e-19
cc_47 N_VDD_c_15_p N_VSS_c_187_n 0.003995f
cc_48 N_VDD_c_48_p N_VSS_c_187_n 0.00163298f
cc_49 N_VDD_c_12_p N_VSS_c_189_n 0.00401122f
cc_50 N_VDD_c_3_p N_VSS_c_189_n 0.0013091f
cc_51 N_VDD_c_51_p N_VSS_c_189_n 0.0010079f
cc_52 N_VDD_c_12_p N_VSS_c_192_n 0.00176255f
cc_53 N_VDD_c_15_p N_VSS_c_193_n 0.00131941f
cc_54 N_VDD_c_16_p N_VSS_c_193_n 0.00593836f
cc_55 N_VDD_c_55_p N_VSS_c_193_n 0.00111239f
cc_56 N_VDD_c_3_p N_VSS_c_196_n 0.0013091f
cc_57 N_VDD_c_8_p N_VSS_c_196_n 0.00841532f
cc_58 N_VDD_c_58_p N_VSS_c_196_n 9.6871e-19
cc_59 N_VDD_c_16_p N_VSS_c_199_n 0.00454933f
cc_60 N_VDD_c_34_p N_VSS_c_200_n 5.34009e-19
cc_61 N_VDD_c_9_p N_VSS_c_201_n 0.00304617f
cc_62 N_VDD_c_6_p N_VSS_c_202_n 2.5062e-19
cc_63 N_VDD_c_9_p N_VSS_c_202_n 0.00529507f
cc_64 N_VDD_c_32_p N_VSS_c_202_n 0.00267625f
cc_65 N_VDD_c_65_p N_VSS_c_202_n 0.0010706f
cc_66 N_VDD_c_15_p N_VSS_c_206_n 7.74609e-19
cc_67 N_VDD_c_3_p N_VSS_c_207_n 0.00104966f
cc_68 N_VDD_c_16_p N_VSS_c_208_n 7.61747e-19
cc_69 N_VDD_c_9_p N_VSS_c_209_n 8.91588e-19
cc_70 N_VDD_c_21_p N_ZI_XI6.X0_CG 9.92565e-19
cc_71 N_VDD_XI2.X0_S N_ZI_XI3.X0_D 3.43419e-19
cc_72 N_VDD_XI0.X0_S N_ZI_XI3.X0_D 3.43419e-19
cc_73 N_VDD_c_6_p N_ZI_XI3.X0_D 3.48267e-19
cc_74 N_VDD_c_34_p N_ZI_XI3.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_PGD N_ZI_c_278_n 2.22031e-19
cc_76 N_VDD_XI6.X0_PGD N_ZI_c_278_n 3.91104e-19
cc_77 N_VDD_c_8_p N_ZI_c_280_n 5.01863e-19
cc_78 N_VDD_c_9_p N_ZI_c_280_n 4.66891e-19
cc_79 N_VDD_XI2.X0_S N_ZI_c_282_n 3.48267e-19
cc_80 N_VDD_XI0.X0_S N_ZI_c_282_n 3.48267e-19
cc_81 N_VDD_c_6_p N_ZI_c_282_n 4.97272e-19
cc_82 N_VDD_c_16_p N_ZI_c_282_n 5.01863e-19
cc_83 N_VDD_c_34_p N_ZI_c_282_n 5.226e-19
cc_84 N_VDD_c_25_p N_ZI_c_287_n 5.3845e-19
cc_85 N_VDD_c_15_p N_ZI_c_288_n 3.65425e-19
cc_86 N_VDD_XI7.X0_D N_Z_XI7.X0_S 3.43419e-19
cc_87 N_VDD_c_12_p N_Z_XI7.X0_S 3.7884e-19
cc_88 N_VDD_c_17_p N_Z_XI7.X0_S 3.72199e-19
cc_89 N_VDD_XI7.X0_D Z 3.48267e-19
cc_90 N_VDD_c_12_p Z 5.12447e-19
cc_91 N_VDD_c_17_p Z 7.4527e-19
cc_92 N_VDD_XI2.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_93 N_VDD_c_15_p N_SELI_XI1.X0_D 3.7884e-19
cc_94 N_VDD_c_6_p N_SELI_XI1.X0_D 3.48267e-19
cc_95 N_VDD_c_95_p N_SELI_XI5.X0_CG 0.00237871f
cc_96 N_VDD_XI2.X0_S N_SELI_c_356_n 3.48267e-19
cc_97 N_VDD_c_15_p N_SELI_c_356_n 5.34458e-19
cc_98 N_VDD_c_6_p N_SELI_c_356_n 6.883e-19
cc_99 N_VDD_XI6.X0_PGD N_SELI_c_359_n 2.27908e-19
cc_100 N_VDD_c_15_p N_SELI_c_359_n 2.61043e-19
cc_101 N_VDD_c_20_p N_SELI_c_359_n 5.3241e-19
cc_102 N_VDD_c_3_p N_SELI_c_359_n 2.36369e-19
cc_103 N_VDD_c_21_p N_SELI_c_359_n 3.99122e-19
cc_104 N_VDD_c_9_p N_SELI_c_364_n 4.30008e-19
cc_105 N_VDD_c_28_p N_SELI_c_365_n 7.54639e-19
cc_106 N_VDD_c_95_p N_SELI_c_365_n 5.0614e-19
cc_107 N_VDD_c_28_p N_SELI_c_367_n 4.85469e-19
cc_108 N_VDD_c_95_p N_SELI_c_367_n 0.0014909f
cc_109 N_VDD_c_25_p N_SEL_XI1.X0_CG 9.92565e-19
cc_110 N_VDD_XI1.X0_PGD N_SEL_c_434_n 4.04053e-19
cc_111 N_VDD_XI6.X0_PGD N_SEL_c_434_n 2.07349e-19
cc_112 N_VDD_XI2.X0_S N_SEL_c_436_n 9.18655e-19
cc_113 N_VDD_c_6_p N_SEL_c_436_n 0.00151457f
cc_114 N_VDD_c_16_p N_SEL_c_438_n 4.35337e-19
cc_115 N_VDD_c_9_p N_SEL_c_439_n 4.25334e-19
cc_116 N_VDD_c_16_p N_SEL_c_440_n 2.49768e-19
cc_117 N_VDD_c_8_p N_SEL_c_440_n 4.35337e-19
cc_118 N_VDD_c_9_p N_SEL_c_442_n 8.17234e-19
cc_119 N_VDD_c_21_p N_SEL_c_443_n 4.93609e-19
cc_120 N_VDD_c_95_p N_SEL_c_444_n 2.00604e-19
cc_121 N_VDD_XI4.X0_PGD N_SEL_c_445_n 3.11814e-19
cc_122 N_VDD_c_9_p N_SEL_c_445_n 3.66936e-19
cc_123 N_VDD_c_6_p N_B_XI5.X0_PGS 2.48132e-19
cc_124 N_VDD_c_6_p B 0.0014278f
cc_125 N_VDD_c_16_p B 0.00141439f
cc_126 N_VDD_c_6_p N_B_c_514_n 9.67317e-19
cc_127 N_VDD_c_16_p N_B_c_514_n 0.00117371f
cc_128 N_VDD_XI4.X0_PGD N_A_XI4.X0_PGS 0.00162178f
cc_129 N_VDD_c_9_p N_A_XI4.X0_PGS 9.35727e-19
cc_130 N_VDD_c_8_p N_A_c_544_n 3.3974e-19
cc_131 N_VDD_c_9_p N_A_c_544_n 4.15738e-19
cc_132 N_VDD_c_28_p A 5.43314e-19
cc_133 N_VDD_c_8_p A 0.00141439f
cc_134 N_VDD_c_9_p A 5.30212e-19
cc_135 N_VDD_c_95_p A 3.48267e-19
cc_136 N_VDD_c_136_p N_A_c_550_n 0.00480616f
cc_137 N_VDD_c_28_p N_A_c_550_n 4.04186e-19
cc_138 N_VDD_c_8_p N_A_c_550_n 0.00117371f
cc_139 N_VDD_c_9_p N_A_c_550_n 3.66936e-19
cc_140 N_VDD_c_95_p N_A_c_550_n 6.39485e-19
cc_141 N_VSS_c_176_n N_ZI_XI7.X0_CG 0.00234241f
cc_142 N_VSS_XI6.X0_S N_ZI_XI5.X0_D 3.43419e-19
cc_143 N_VSS_XI4.X0_S N_ZI_XI5.X0_D 3.43419e-19
cc_144 N_VSS_c_173_n N_ZI_XI5.X0_D 3.48267e-19
cc_145 N_VSS_XI7.X0_PGS N_ZI_c_278_n 3.99472e-19
cc_146 N_VSS_c_158_n N_ZI_c_294_n 0.00126951f
cc_147 N_VSS_c_176_n N_ZI_c_294_n 8.72558e-19
cc_148 N_VSS_XI6.X0_S N_ZI_c_280_n 3.48267e-19
cc_149 N_VSS_XI4.X0_S N_ZI_c_280_n 3.48267e-19
cc_150 N_VSS_c_166_n N_ZI_c_280_n 0.00100597f
cc_151 N_VSS_c_173_n N_ZI_c_280_n 4.40384e-19
cc_152 N_VSS_c_196_n N_ZI_c_280_n 5.12922e-19
cc_153 N_VSS_c_200_n N_ZI_c_280_n 6.1924e-19
cc_154 N_VSS_c_202_n N_ZI_c_280_n 0.00113121f
cc_155 N_VSS_c_193_n N_ZI_c_282_n 5.12922e-19
cc_156 N_VSS_c_158_n N_ZI_c_287_n 4.56568e-19
cc_157 N_VSS_c_176_n N_ZI_c_287_n 0.0014909f
cc_158 N_VSS_c_162_n N_ZI_c_288_n 4.17431e-19
cc_159 N_VSS_c_166_n N_ZI_c_288_n 6.40656e-19
cc_160 N_VSS_c_189_n N_ZI_c_288_n 0.00101727f
cc_161 N_VSS_c_193_n N_ZI_c_288_n 0.00147997f
cc_162 N_VSS_c_196_n N_ZI_c_288_n 2.59546e-19
cc_163 N_VSS_c_187_n N_ZI_c_311_n 0.0011789f
cc_164 N_VSS_XI6.X0_S N_Z_XI7.X0_S 3.43419e-19
cc_165 N_VSS_c_166_n N_Z_XI7.X0_S 3.48267e-19
cc_166 N_VSS_XI6.X0_S Z 3.48267e-19
cc_167 N_VSS_c_166_n Z 7.85754e-19
cc_168 N_VSS_XI1.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_169 N_VSS_c_157_n N_SELI_XI1.X0_D 3.48267e-19
cc_170 N_VSS_c_184_n N_SELI_c_371_n 0.00234241f
cc_171 N_VSS_c_157_n N_SELI_c_356_n 6.0686e-19
cc_172 N_VSS_c_166_n N_SELI_c_359_n 0.00130595f
cc_173 N_VSS_c_189_n N_SELI_c_359_n 4.10258e-19
cc_174 N_VSS_c_170_n N_SELI_c_364_n 0.00135778f
cc_175 N_VSS_c_184_n N_SELI_c_364_n 4.99367e-19
cc_176 N_VSS_c_196_n N_SELI_c_364_n 4.69529e-19
cc_177 N_VSS_c_202_n N_SELI_c_364_n 9.62347e-19
cc_178 N_VSS_c_170_n N_SELI_c_379_n 4.56568e-19
cc_179 N_VSS_c_184_n N_SELI_c_379_n 0.0014909f
cc_180 N_VSS_c_196_n N_SELI_c_381_n 7.6099e-19
cc_181 N_VSS_c_202_n N_SELI_c_381_n 6.2582e-19
cc_182 N_VSS_XI7.X0_PGS N_SEL_c_434_n 2.22031e-19
cc_183 N_VSS_XI2.X0_PGD N_SEL_c_434_n 3.91879e-19
cc_184 N_VSS_c_180_n N_SEL_c_449_n 0.00272336f
cc_185 N_VSS_c_193_n N_SEL_c_436_n 4.08267e-19
cc_186 N_VSS_c_202_n N_SEL_c_439_n 2.03139e-19
cc_187 N_VSS_c_196_n N_SEL_c_440_n 2.53418e-19
cc_188 N_VSS_c_257_p N_SEL_c_453_n 3.73191e-19
cc_189 N_VSS_c_162_n N_SEL_c_453_n 6.21258e-19
cc_190 N_VSS_c_162_n N_SEL_c_443_n 4.56568e-19
cc_191 N_VSS_c_180_n N_SEL_c_443_n 0.0014909f
cc_192 N_VSS_XI3.X0_PGD N_SEL_c_444_n 3.11814e-19
cc_193 N_VSS_c_184_n N_SEL_c_445_n 2.00604e-19
cc_194 N_VSS_XI2.X0_PGS N_B_XI5.X0_PGS 0.00172969f
cc_195 N_VSS_XI3.X0_PGD N_B_XI5.X0_PGS 0.00152606f
cc_196 N_VSS_c_265_p N_B_c_518_n 0.00172969f
cc_197 N_VSS_c_170_n B 3.98896e-19
cc_198 N_VSS_c_184_n B 3.5189e-19
cc_199 N_VSS_c_156_n N_B_c_514_n 0.00295829f
cc_200 N_VSS_c_170_n N_B_c_514_n 3.5189e-19
cc_201 N_VSS_c_180_n N_B_c_514_n 7.89771e-19
cc_202 N_VSS_c_184_n N_B_c_514_n 6.80896e-19
cc_203 N_VSS_c_196_n A 2.11858e-19
cc_204 N_ZI_c_282_n N_SELI_c_356_n 3.26181e-19
cc_205 N_ZI_c_288_n N_SELI_c_356_n 0.00213954f
cc_206 N_ZI_c_278_n N_SELI_c_359_n 4.92356e-19
cc_207 N_ZI_c_288_n N_SELI_c_359_n 0.00182433f
cc_208 N_ZI_c_278_n N_SELI_c_387_n 2.38253e-19
cc_209 N_ZI_c_294_n N_SELI_c_387_n 0.00150231f
cc_210 N_ZI_c_287_n N_SELI_c_387_n 0.00110082f
cc_211 N_ZI_c_282_n N_SELI_c_364_n 0.00173524f
cc_212 N_ZI_c_280_n N_SELI_c_365_n 0.00183505f
cc_213 N_ZI_c_288_n N_SELI_c_365_n 0.00144518f
cc_214 N_ZI_c_280_n N_SELI_c_381_n 7.38292e-19
cc_215 N_ZI_c_288_n N_SELI_c_381_n 7.7914e-19
cc_216 N_ZI_c_280_n N_SELI_c_395_n 5.82645e-19
cc_217 N_ZI_c_282_n N_SELI_c_395_n 3.22755e-19
cc_218 N_ZI_c_326_p N_SELI_c_395_n 6.45182e-19
cc_219 N_ZI_c_282_n N_SELI_c_398_n 7.64986e-19
cc_220 N_ZI_c_278_n N_SEL_c_434_n 0.00371647f
cc_221 N_ZI_c_287_n N_SEL_c_460_n 3.81736e-19
cc_222 N_ZI_XI3.X0_D N_SEL_c_438_n 9.94581e-19
cc_223 N_ZI_c_282_n N_SEL_c_438_n 0.00247421f
cc_224 N_ZI_c_280_n N_SEL_c_439_n 6.15647e-19
cc_225 N_ZI_c_326_p N_SEL_c_439_n 0.00107464f
cc_226 N_ZI_XI5.X0_D N_SEL_c_465_n 9.94581e-19
cc_227 N_ZI_c_280_n N_SEL_c_465_n 0.00243387f
cc_228 N_ZI_c_288_n N_SEL_c_453_n 0.00217047f
cc_229 N_ZI_c_282_n N_SEL_c_468_n 2.25033e-19
cc_230 N_ZI_c_278_n N_SEL_c_443_n 3.81736e-19
cc_231 N_ZI_XI6.X0_CG N_B_XI5.X0_PGS 0.00182649f
cc_232 N_Z_XI7.X0_S N_SELI_c_387_n 9.09799e-19
cc_233 Z N_SELI_c_387_n 0.00147087f
cc_234 N_SELI_c_356_n N_SEL_c_434_n 8.51271e-19
cc_235 N_SELI_c_365_n N_SEL_c_436_n 0.00269197f
cc_236 N_SELI_c_364_n N_SEL_c_438_n 0.00117605f
cc_237 N_SELI_c_356_n N_SEL_c_439_n 2.52418e-19
cc_238 N_SELI_c_364_n N_SEL_c_440_n 3.73414e-19
cc_239 N_SELI_c_365_n N_SEL_c_465_n 0.00160262f
cc_240 N_SELI_c_367_n N_SEL_c_465_n 9.78333e-19
cc_241 N_SELI_c_356_n N_SEL_c_453_n 0.00246582f
cc_242 N_SELI_c_359_n N_SEL_c_453_n 0.00269197f
cc_243 N_SELI_c_364_n N_SEL_c_468_n 2.32653e-19
cc_244 N_SELI_c_379_n N_SEL_c_468_n 3.48267e-19
cc_245 N_SELI_c_364_n N_SEL_c_442_n 9.4965e-19
cc_246 N_SELI_c_365_n N_SEL_c_442_n 2.32653e-19
cc_247 N_SELI_c_367_n N_SEL_c_442_n 3.48267e-19
cc_248 N_SELI_c_356_n N_SEL_c_443_n 9.71051e-19
cc_249 N_SELI_c_359_n N_SEL_c_443_n 6.26941e-19
cc_250 N_SELI_c_364_n N_SEL_c_444_n 3.48267e-19
cc_251 N_SELI_c_365_n N_SEL_c_444_n 7.22902e-19
cc_252 N_SELI_c_367_n N_SEL_c_444_n 0.0049864f
cc_253 N_SELI_c_379_n N_SEL_c_444_n 9.11855e-19
cc_254 N_SELI_c_364_n N_SEL_c_445_n 4.99367e-19
cc_255 N_SELI_c_365_n N_SEL_c_445_n 3.68647e-19
cc_256 N_SELI_c_367_n N_SEL_c_445_n 9.28301e-19
cc_257 N_SELI_c_379_n N_SEL_c_445_n 0.00490516f
cc_258 N_SELI_XI5.X0_CG N_B_XI5.X0_PGS 4.41254e-19
cc_259 N_SELI_c_356_n N_B_XI5.X0_PGS 2.21243e-19
cc_260 N_SELI_c_359_n N_B_XI5.X0_PGS 7.89402e-19
cc_261 N_SELI_c_367_n N_B_XI5.X0_PGS 0.00186882f
cc_262 N_SELI_c_367_n N_B_c_514_n 2.00604e-19
cc_263 N_SELI_c_371_n N_A_XI4.X0_PGS 4.65768e-19
cc_264 N_SELI_c_379_n N_A_XI4.X0_PGS 0.00276355f
cc_265 N_SELI_c_379_n N_A_c_550_n 2.00604e-19
cc_266 N_SEL_c_449_n N_B_XI5.X0_PGS 2.07014e-19
cc_267 N_SEL_c_495_p N_B_XI5.X0_PGS 4.3669e-19
cc_268 N_SEL_c_436_n N_B_XI5.X0_PGS 7.4877e-19
cc_269 N_SEL_c_443_n N_B_XI5.X0_PGS 0.00100354f
cc_270 N_SEL_c_444_n N_B_XI5.X0_PGS 0.00202689f
cc_271 N_SEL_c_468_n B 6.87706e-19
cc_272 N_SEL_c_444_n B 4.56568e-19
cc_273 N_SEL_c_495_p N_B_c_514_n 0.00234241f
cc_274 N_SEL_c_468_n N_B_c_514_n 5.02946e-19
cc_275 N_SEL_c_444_n N_B_c_514_n 0.0014909f
cc_276 N_SEL_XI4.X0_CG N_A_XI4.X0_PGS 4.54863e-19
cc_277 N_SEL_c_445_n N_A_XI4.X0_PGS 0.00276355f
cc_278 N_SEL_c_442_n A 7.05846e-19
cc_279 N_SEL_c_445_n A 4.56568e-19
cc_280 N_SEL_XI4.X0_CG N_A_c_550_n 0.00234241f
cc_281 N_SEL_c_442_n N_A_c_550_n 5.02946e-19
cc_282 N_SEL_c_445_n N_A_c_550_n 0.0014909f
cc_283 N_B_XI5.X0_PGS N_A_XI4.X0_PGS 0.00137635f
*
.ends
*
*
.subckt MUX2_HPNW4 A B S0 Y VDD VSS
xgate (VDD VSS Y S0 B A) G4_MUX2_N1
.ends
*
* File: G3_MUXI2_N1.pex.netlist
* Created: Wed Mar  9 13:36:32 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MUXI2_N1_VSS 2 4 6 8 10 12 14 29 31 39 63 68 73 78 83 92 101 110
+ 115 121 127 133 135 140 142 144 145 146 147 Vss
c86 147 Vss 4.28045e-19
c87 146 Vss 3.62111e-19
c88 145 Vss 3.75522e-19
c89 142 Vss 0.00430383f
c90 140 Vss 0.00143623f
c91 135 Vss 0.00139741f
c92 133 Vss 0.002505f
c93 128 Vss 0.00127887f
c94 127 Vss 0.00644124f
c95 121 Vss 0.00399642f
c96 116 Vss 0.0013489f
c97 115 Vss 0.00539877f
c98 110 Vss 0.00225019f
c99 109 Vss 0.00129191f
c100 101 Vss 0.00660977f
c101 92 Vss 0.00400552f
c102 83 Vss 1.70165e-19
c103 78 Vss 0.00106984f
c104 73 Vss 0.00241148f
c105 68 Vss 2.9197e-19
c106 63 Vss 0.00126608f
c107 45 Vss 0.0785271f
c108 39 Vss 0.0343198f
c109 38 Vss 0.0688517f
c110 31 Vss 7.82991e-20
c111 29 Vss 0.0338093f
c112 28 Vss 0.0998552f
c113 14 Vss 0.0835744f
c114 12 Vss 0.00226958f
c115 10 Vss 0.0837985f
c116 8 Vss 7.32238e-19
c117 6 Vss 0.0838866f
c118 4 Vss 0.0825199f
c119 2 Vss 0.00266844f
r120 141 147 0.551426
r121 141 142 13.3371
r122 140 147 0.551426
r123 139 140 4.16786
r124 135 147 0.0828784
r125 134 146 0.494161
r126 133 142 0.652036
r127 133 134 4.41793
r128 129 146 0.128424
r129 127 139 0.652036
r130 127 128 13.0037
r131 123 128 0.652036
r132 122 145 0.494161
r133 121 146 0.494161
r134 121 122 10.2946
r135 117 145 0.128424
r136 115 145 0.494161
r137 115 116 10.1279
r138 111 144 0.306046
r139 110 116 0.652036
r140 109 144 0.349767
r141 109 110 4.16786
r142 83 135 1.82344
r143 78 101 1.16709
r144 78 129 2.16729
r145 73 123 4.83471
r146 68 92 1.16709
r147 68 117 2.16729
r148 63 111 1.82344
r149 45 101 0.238214
r150 43 45 1.8672
r151 40 43 0.0685365
r152 38 43 0.5835
r153 38 39 2.8008
r154 35 39 0.652036
r155 31 92 0.238214
r156 29 31 1.45875
r157 28 32 0.652036
r158 28 31 1.45875
r159 25 29 0.652036
r160 14 40 2.5674
r161 12 83 1.16709
r162 10 35 2.5674
r163 8 73 1.16709
r164 6 32 2.5674
r165 4 25 2.5674
r166 2 63 1.16709
.ends

.subckt PM_G3_MUXI2_N1_VDD 2 4 6 8 12 14 28 38 60 62 63 66 68 72 74 75 76 77 78
+ 79 81 82 87 88 90 99 Vss
c99 99 Vss 0.00651319f
c100 90 Vss 0.00555165f
c101 88 Vss 3.54369e-19
c102 82 Vss 4.42156e-19
c103 81 Vss 0.00190072f
c104 79 Vss 0.00690705f
c105 78 Vss 8.63529e-19
c106 77 Vss 4.40622e-19
c107 76 Vss 0.00130949f
c108 75 Vss 6.09322e-19
c109 74 Vss 0.00547771f
c110 72 Vss 9.38425e-19
c111 68 Vss 0.00834424f
c112 66 Vss 0.00132511f
c113 63 Vss 6.1175e-19
c114 62 Vss 0.00344974f
c115 60 Vss 0.00121763f
c116 39 Vss 0.0805612f
c117 38 Vss 0.102888f
c118 29 Vss 0.0355046f
c119 28 Vss 0.1003f
c120 14 Vss 0.00271849f
c121 12 Vss 0.0806222f
c122 8 Vss 0.0814405f
c123 6 Vss 0.00155055f
c124 4 Vss 0.0842982f
c125 2 Vss 0.0825186f
r126 80 88 0.537385
r127 80 81 4.16786
r128 79 88 0.537385
r129 78 87 0.326018
r130 78 79 13.3788
r131 77 84 0.510562
r132 76 88 0.0936215
r133 76 77 1.35523
r134 74 87 0.326018
r135 74 75 10.1279
r136 72 99 1.16709
r137 70 75 0.652036
r138 70 72 2.16729
r139 69 82 0.494161
r140 68 81 0.652036
r141 68 69 13.0037
r142 64 82 0.128424
r143 64 66 4.83471
r144 62 82 0.494161
r145 62 63 7.46046
r146 60 90 1.16709
r147 58 63 0.652036
r148 58 60 2.16729
r149 44 99 0.238214
r150 44 46 1.92555
r151 39 46 0.5835
r152 38 40 0.652036
r153 38 39 2.8008
r154 35 46 0.0685365
r155 31 90 0.238214
r156 29 31 1.45875
r157 28 32 0.652036
r158 28 31 1.45875
r159 25 29 0.652036
r160 14 84 1.16709
r161 12 40 2.5674
r162 8 35 2.5674
r163 6 66 1.16709
r164 4 25 2.5674
r165 2 32 2.5674
.ends

.subckt PM_G3_MUXI2_N1_SELI 2 6 8 21 33 35 38 43 53 58 72 77 78 Vss
c67 78 Vss 3.71671e-19
c68 72 Vss 0.00114167f
c69 58 Vss 0.00216403f
c70 53 Vss 0.00206075f
c71 43 Vss 9.19217e-19
c72 38 Vss 0.00147194f
c73 36 Vss 0.00160147f
c74 35 Vss 0.00416276f
c75 33 Vss 0.00272744f
c76 21 Vss 0.0575023f
c77 6 Vss 0.0575023f
c78 2 Vss 0.00148239f
r79 77 78 0.655813
r80 76 77 3.501
r81 72 76 0.655813
r82 43 53 1.16709
r83 43 72 2.00578
r84 43 46 0.833571
r85 38 58 1.16709
r86 38 78 2.00578
r87 35 46 0.0685365
r88 35 36 7.46046
r89 31 36 0.652036
r90 31 33 5.58493
r91 21 58 0.50025
r92 18 53 0.50025
r93 8 21 1.80885
r94 6 18 1.80885
r95 2 33 1.16709
.ends

.subckt PM_G3_MUXI2_N1_SEL 2 4 6 8 16 22 26 36 37 40 42 46 51 58 63 68 72 77 78
+ Vss
c73 78 Vss 8.48303e-20
c74 77 Vss 2.4421e-20
c75 72 Vss 7.30413e-19
c76 68 Vss 0.00150427f
c77 63 Vss 0.00289461f
c78 58 Vss 0.00236419f
c79 51 Vss 4.10742e-19
c80 46 Vss 1.61132e-19
c81 42 Vss 0.00131501f
c82 37 Vss 0.00193143f
c83 36 Vss 6.68718e-20
c84 26 Vss 0.057622f
c85 22 Vss 0.0712295f
c86 20 Vss 0.0247918f
c87 17 Vss 0.0369263f
c88 16 Vss 0.187844f
c89 8 Vss 0.0575023f
c90 2 Vss 0.084915f
r91 76 78 0.655813
r92 76 77 3.501
r93 72 77 0.655813
r94 54 63 1.16709
r95 54 72 2.00578
r96 51 54 0.5835
r97 49 58 1.16709
r98 46 49 0.5835
r99 42 68 1.16709
r100 42 78 2.00578
r101 38 46 0.0685365
r102 38 40 1.70882
r103 37 51 0.0685365
r104 37 40 2.87582
r105 36 58 0.0476429
r106 33 68 0.50025
r107 26 63 0.50025
r108 22 58 0.357321
r109 20 36 0.326018
r110 20 22 0.40845
r111 17 36 6.7686
r112 16 36 0.326018
r113 16 36 0.1167
r114 13 17 0.652036
r115 8 33 1.80885
r116 6 26 1.80885
r117 4 22 2.15895
r118 2 13 2.5674
.ends

.subckt PM_G3_MUXI2_N1_B 2 4 7 16 20 24 27 Vss
c22 27 Vss 0.00591505f
c23 24 Vss 5.28389e-19
c24 20 Vss 0.0298499f
c25 16 Vss 0.0664813f
c26 7 Vss 0.142354f
c27 4 Vss 0.272228f
c28 2 Vss 0.0800936f
r29 24 27 1.16709
r30 16 27 0.50025
r31 16 18 1.9839
r32 12 20 0.494161
r33 9 20 0.494161
r34 8 18 0.0685365
r35 7 20 0.128424
r36 7 8 4.7847
r37 4 12 9.04425
r38 2 9 2.62575
.ends

.subckt PM_G3_MUXI2_N1_Z 2 4 30 33 Vss
c33 30 Vss 0.00283949f
c34 4 Vss 0.00148239f
c35 2 Vss 0.00156677f
r36 33 35 5.16814
r37 30 33 4.00114
r38 4 35 1.16709
r39 2 30 1.16709
.ends

.subckt PM_G3_MUXI2_N1_A 2 4 14 19 22 Vss
c24 22 Vss 0.00548526f
c25 19 Vss 4.55558e-19
c26 14 Vss 0.0830192f
c27 2 Vss 0.4453f
r28 19 22 1.16709
r29 12 22 0.238214
r30 12 14 1.92555
r31 7 14 0.0685365
r32 2 4 12.837
r33 2 7 2.5674
.ends

.subckt G3_MUXI2_N1  VSS VDD SEL B Z A
*
* A	A
* Z	Z
* B	B
* SEL	SEL
* VDD	VDD
* VSS	VSS
XI1.X0 N_SELI_XI1.X0_D N_VDD_XI1.X0_PGD N_SEL_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI2.X0 N_SELI_XI1.X0_D N_VSS_XI2.X0_PGD N_SEL_XI2.X0_CG N_VSS_XI2.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_SELI_XI5.X0_CG N_B_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW4
XI3.X0 N_Z_XI3.X0_D N_VSS_XI3.X0_PGD N_SEL_XI3.X0_CG N_B_XI3.X0_PGS
+ N_VDD_XI2.X0_S TIGFET_HPNW4
XI4.X0 N_Z_XI5.X0_D N_VDD_XI4.X0_PGD N_SEL_XI4.X0_CG N_A_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW4
XI0.X0 N_Z_XI3.X0_D N_VSS_XI0.X0_PGD N_SELI_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW4
*
x_PM_G3_MUXI2_N1_VSS N_VSS_XI1.X0_S N_VSS_XI2.X0_PGD N_VSS_XI2.X0_PGS
+ N_VSS_XI5.X0_S N_VSS_XI3.X0_PGD N_VSS_XI4.X0_S N_VSS_XI0.X0_PGD N_VSS_c_4_p
+ N_VSS_c_62_p N_VSS_c_21_p N_VSS_c_47_p N_VSS_c_5_p N_VSS_c_27_p N_VSS_c_18_p
+ N_VSS_c_29_p N_VSS_c_6_p N_VSS_c_20_p N_VSS_c_7_p N_VSS_c_11_p N_VSS_c_12_p
+ N_VSS_c_30_p N_VSS_c_25_p N_VSS_c_32_p N_VSS_c_37_p N_VSS_c_38_p VSS
+ N_VSS_c_13_p N_VSS_c_26_p N_VSS_c_39_p Vss PM_G3_MUXI2_N1_VSS
x_PM_G3_MUXI2_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI2.X0_S
+ N_VDD_XI5.X0_PGD N_VDD_XI4.X0_PGD N_VDD_XI0.X0_S N_VDD_c_90_n N_VDD_c_181_p
+ N_VDD_c_91_n N_VDD_c_94_n N_VDD_c_100_n N_VDD_c_101_n N_VDD_c_107_n
+ N_VDD_c_113_n N_VDD_c_114_n N_VDD_c_117_n N_VDD_c_118_n N_VDD_c_119_n
+ N_VDD_c_120_n N_VDD_c_121_n N_VDD_c_126_n N_VDD_c_128_n VDD N_VDD_c_129_n
+ N_VDD_c_130_n N_VDD_c_135_p Vss PM_G3_MUXI2_N1_VDD
x_PM_G3_MUXI2_N1_SELI N_SELI_XI1.X0_D N_SELI_XI5.X0_CG N_SELI_XI0.X0_CG
+ N_SELI_c_188_n N_SELI_c_189_n N_SELI_c_192_n N_SELI_c_193_n N_SELI_c_209_n
+ N_SELI_c_211_n N_SELI_c_196_n N_SELI_c_198_n N_SELI_c_199_n N_SELI_c_231_p Vss
+ PM_G3_MUXI2_N1_SELI
x_PM_G3_MUXI2_N1_SEL N_SEL_XI1.X0_CG N_SEL_XI2.X0_CG N_SEL_XI3.X0_CG
+ N_SEL_XI4.X0_CG N_SEL_c_253_n N_SEL_c_254_n N_SEL_c_305_p N_SEL_c_255_n
+ N_SEL_c_257_n SEL N_SEL_c_258_n N_SEL_c_259_n N_SEL_c_274_n N_SEL_c_260_n
+ N_SEL_c_275_n N_SEL_c_262_n N_SEL_c_263_n N_SEL_c_265_n N_SEL_c_266_n Vss
+ PM_G3_MUXI2_N1_SEL
x_PM_G3_MUXI2_N1_B N_B_XI5.X0_PGS N_B_XI3.X0_PGS N_B_c_326_n N_B_c_344_n
+ N_B_c_336_n B N_B_c_328_n Vss PM_G3_MUXI2_N1_B
x_PM_G3_MUXI2_N1_Z N_Z_XI5.X0_D N_Z_XI3.X0_D N_Z_c_352_n Z Vss PM_G3_MUXI2_N1_Z
x_PM_G3_MUXI2_N1_A N_A_XI4.X0_PGS N_A_XI0.X0_PGS N_A_c_383_n A N_A_c_389_n Vss
+ PM_G3_MUXI2_N1_A
cc_1 N_VSS_XI2.X0_PGD N_VDD_XI1.X0_PGD 0.0017188f
cc_2 N_VSS_XI3.X0_PGD N_VDD_XI5.X0_PGD 2.27468e-19
cc_3 N_VSS_XI0.X0_PGD N_VDD_XI4.X0_PGD 2.27468e-19
cc_4 N_VSS_c_4_p N_VDD_c_90_n 0.0017188f
cc_5 N_VSS_c_5_p N_VDD_c_91_n 9.32947e-19
cc_6 N_VSS_c_6_p N_VDD_c_91_n 3.82294e-19
cc_7 N_VSS_c_7_p N_VDD_c_91_n 4.10707e-19
cc_8 N_VSS_c_4_p N_VDD_c_94_n 2.72324e-19
cc_9 N_VSS_c_5_p N_VDD_c_94_n 0.00141228f
cc_10 N_VSS_c_6_p N_VDD_c_94_n 0.00112249f
cc_11 N_VSS_c_11_p N_VDD_c_94_n 0.00419135f
cc_12 N_VSS_c_12_p N_VDD_c_94_n 0.00124457f
cc_13 N_VSS_c_13_p N_VDD_c_94_n 7.74609e-19
cc_14 N_VSS_c_11_p N_VDD_c_100_n 0.00157719f
cc_15 N_VSS_XI2.X0_PGS N_VDD_c_101_n 2.93604e-19
cc_16 N_VSS_XI3.X0_PGD N_VDD_c_101_n 2.36238e-19
cc_17 N_VSS_c_5_p N_VDD_c_101_n 0.00181129f
cc_18 N_VSS_c_18_p N_VDD_c_101_n 7.45025e-19
cc_19 N_VSS_c_6_p N_VDD_c_101_n 9.55109e-19
cc_20 N_VSS_c_20_p N_VDD_c_101_n 2.60394e-19
cc_21 N_VSS_c_21_p N_VDD_c_107_n 0.00102426f
cc_22 N_VSS_c_18_p N_VDD_c_107_n 0.00161703f
cc_23 N_VSS_c_20_p N_VDD_c_107_n 2.03837e-19
cc_24 N_VSS_c_12_p N_VDD_c_107_n 0.0056811f
cc_25 N_VSS_c_25_p N_VDD_c_107_n 0.00454933f
cc_26 N_VSS_c_26_p N_VDD_c_107_n 7.61747e-19
cc_27 N_VSS_c_27_p N_VDD_c_113_n 0.00125492f
cc_28 N_VSS_XI4.X0_S N_VDD_c_114_n 3.7884e-19
cc_29 N_VSS_c_29_p N_VDD_c_114_n 4.73473e-19
cc_30 N_VSS_c_30_p N_VDD_c_114_n 0.00742779f
cc_31 N_VSS_c_30_p N_VDD_c_117_n 0.00149994f
cc_32 N_VSS_c_32_p N_VDD_c_118_n 4.31398e-19
cc_33 N_VSS_c_29_p N_VDD_c_119_n 2.14355e-19
cc_34 N_VSS_c_30_p N_VDD_c_120_n 0.00106317f
cc_35 N_VSS_XI4.X0_S N_VDD_c_121_n 9.5668e-19
cc_36 N_VSS_c_29_p N_VDD_c_121_n 0.00165395f
cc_37 N_VSS_c_37_p N_VDD_c_121_n 0.00364836f
cc_38 N_VSS_c_38_p N_VDD_c_121_n 0.0050309f
cc_39 N_VSS_c_39_p N_VDD_c_121_n 8.91588e-19
cc_40 N_VSS_c_18_p N_VDD_c_126_n 4.6996e-19
cc_41 N_VSS_c_38_p N_VDD_c_126_n 0.00295094f
cc_42 N_VSS_c_12_p N_VDD_c_128_n 0.00112088f
cc_43 N_VSS_c_38_p N_VDD_c_129_n 9.75645e-19
cc_44 N_VSS_c_5_p N_VDD_c_130_n 3.48267e-19
cc_45 N_VSS_c_6_p N_VDD_c_130_n 8.0279e-19
cc_46 N_VSS_XI1.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_47 N_VSS_c_47_p N_SELI_XI1.X0_D 3.48267e-19
cc_48 N_VSS_c_20_p N_SELI_c_188_n 0.00234241f
cc_49 N_VSS_XI1.X0_S N_SELI_c_189_n 3.48267e-19
cc_50 N_VSS_c_47_p N_SELI_c_189_n 8.47286e-19
cc_51 N_VSS_c_11_p N_SELI_c_189_n 2.65284e-19
cc_52 N_VSS_c_27_p N_SELI_c_192_n 0.00140233f
cc_53 N_VSS_c_18_p N_SELI_c_193_n 0.00135778f
cc_54 N_VSS_c_20_p N_SELI_c_193_n 4.99367e-19
cc_55 N_VSS_c_38_p N_SELI_c_193_n 9.07743e-19
cc_56 N_VSS_c_18_p N_SELI_c_196_n 4.56568e-19
cc_57 N_VSS_c_20_p N_SELI_c_196_n 0.0014909f
cc_58 N_VSS_c_30_p N_SELI_c_198_n 7.53578e-19
cc_59 N_VSS_c_38_p N_SELI_c_199_n 5.03655e-19
cc_60 N_VSS_XI2.X0_PGD N_SEL_c_253_n 4.12362e-19
cc_61 N_VSS_c_6_p N_SEL_c_254_n 0.00234241f
cc_62 N_VSS_c_62_p N_SEL_c_255_n 9.36847e-19
cc_63 N_VSS_c_6_p N_SEL_c_255_n 2.03369e-19
cc_64 N_VSS_c_12_p N_SEL_c_257_n 5.44326e-19
cc_65 N_VSS_c_38_p N_SEL_c_258_n 3.80099e-19
cc_66 N_VSS_c_5_p N_SEL_c_259_n 8.36018e-19
cc_67 N_VSS_c_5_p N_SEL_c_260_n 4.56568e-19
cc_68 N_VSS_c_6_p N_SEL_c_260_n 6.1245e-19
cc_69 N_VSS_c_20_p N_SEL_c_262_n 2.00604e-19
cc_70 N_VSS_c_12_p N_SEL_c_263_n 0.00127961f
cc_71 N_VSS_c_30_p N_SEL_c_263_n 2.81471e-19
cc_72 N_VSS_c_38_p N_SEL_c_265_n 4.36463e-19
cc_73 N_VSS_c_30_p N_SEL_c_266_n 0.00119312f
cc_74 N_VSS_XI2.X0_PGS N_B_c_326_n 2.96367e-19
cc_75 N_VSS_c_27_p B 0.00220388f
cc_76 N_VSS_XI5.X0_S N_B_c_328_n 0.00246958f
cc_77 N_VSS_c_27_p N_B_c_328_n 8.835e-19
cc_78 N_VSS_XI5.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_79 N_VSS_XI4.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_80 N_VSS_c_27_p N_Z_XI5.X0_D 3.48267e-19
cc_81 N_VSS_c_29_p N_Z_XI5.X0_D 3.48267e-19
cc_82 N_VSS_XI5.X0_S N_Z_c_352_n 3.48267e-19
cc_83 N_VSS_XI4.X0_S N_Z_c_352_n 3.48267e-19
cc_84 N_VSS_c_27_p N_Z_c_352_n 5.68449e-19
cc_85 N_VSS_c_29_p N_Z_c_352_n 5.69026e-19
cc_86 N_VSS_c_38_p N_Z_c_352_n 3.26224e-19
cc_87 N_VDD_XI2.X0_S N_SELI_XI1.X0_D 3.43419e-19
cc_88 N_VDD_c_94_n N_SELI_XI1.X0_D 3.7884e-19
cc_89 N_VDD_c_101_n N_SELI_XI1.X0_D 3.48267e-19
cc_90 N_VDD_c_135_p N_SELI_XI5.X0_CG 0.00237871f
cc_91 N_VDD_XI2.X0_S N_SELI_c_189_n 3.48267e-19
cc_92 N_VDD_c_94_n N_SELI_c_189_n 5.34437e-19
cc_93 N_VDD_c_101_n N_SELI_c_189_n 7.03427e-19
cc_94 N_VDD_c_94_n N_SELI_c_192_n 2.96638e-19
cc_95 N_VDD_c_121_n N_SELI_c_193_n 6.15494e-19
cc_96 N_VDD_c_113_n N_SELI_c_209_n 7.54639e-19
cc_97 N_VDD_c_135_p N_SELI_c_209_n 5.0614e-19
cc_98 N_VDD_c_113_n N_SELI_c_211_n 4.85469e-19
cc_99 N_VDD_c_135_p N_SELI_c_211_n 0.013665f
cc_100 N_VDD_c_121_n N_SELI_c_196_n 3.66936e-19
cc_101 N_VDD_c_130_n N_SEL_XI1.X0_CG 8.03148e-19
cc_102 N_VDD_XI1.X0_PGD N_SEL_c_253_n 4.25379e-19
cc_103 N_VDD_XI2.X0_S N_SEL_c_257_n 9.18655e-19
cc_104 N_VDD_c_101_n N_SEL_c_257_n 0.00161606f
cc_105 N_VDD_c_107_n N_SEL_c_258_n 2.90143e-19
cc_106 N_VDD_c_114_n N_SEL_c_258_n 3.06021e-19
cc_107 N_VDD_c_121_n N_SEL_c_258_n 6.68274e-19
cc_108 N_VDD_c_107_n N_SEL_c_274_n 2.1079e-19
cc_109 N_VDD_c_107_n N_SEL_c_275_n 2.19082e-19
cc_110 N_VDD_c_135_p N_SEL_c_275_n 2.00604e-19
cc_111 N_VDD_XI4.X0_PGD N_SEL_c_262_n 3.11814e-19
cc_112 N_VDD_c_121_n N_SEL_c_262_n 3.66936e-19
cc_113 N_VDD_c_107_n N_SEL_c_263_n 4.86613e-19
cc_114 N_VDD_c_121_n N_SEL_c_265_n 2.2501e-19
cc_115 N_VDD_c_114_n N_Z_XI5.X0_D 3.7884e-19
cc_116 N_VDD_XI2.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_117 N_VDD_XI0.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_118 N_VDD_c_101_n N_Z_XI3.X0_D 3.48267e-19
cc_119 N_VDD_c_107_n N_Z_XI3.X0_D 3.7884e-19
cc_120 N_VDD_c_119_n N_Z_XI3.X0_D 3.72199e-19
cc_121 N_VDD_XI2.X0_S N_Z_c_352_n 3.48267e-19
cc_122 N_VDD_XI0.X0_S N_Z_c_352_n 3.48267e-19
cc_123 N_VDD_c_101_n N_Z_c_352_n 8.10024e-19
cc_124 N_VDD_c_107_n N_Z_c_352_n 5.35804e-19
cc_125 N_VDD_c_114_n N_Z_c_352_n 5.35804e-19
cc_126 N_VDD_c_119_n N_Z_c_352_n 8.05266e-19
cc_127 N_VDD_c_121_n N_Z_c_352_n 7.45211e-19
cc_128 N_VDD_XI4.X0_PGD N_A_XI4.X0_PGS 0.00162178f
cc_129 N_VDD_c_121_n N_A_XI4.X0_PGS 0.0010699f
cc_130 N_VDD_c_114_n N_A_c_383_n 3.3974e-19
cc_131 N_VDD_c_121_n N_A_c_383_n 4.15738e-19
cc_132 N_VDD_c_113_n A 5.43314e-19
cc_133 N_VDD_c_114_n A 0.00141439f
cc_134 N_VDD_c_121_n A 5.04211e-19
cc_135 N_VDD_c_135_p A 3.48267e-19
cc_136 N_VDD_c_181_p N_A_c_389_n 0.00480616f
cc_137 N_VDD_c_113_n N_A_c_389_n 3.89161e-19
cc_138 N_VDD_c_114_n N_A_c_389_n 0.00117371f
cc_139 N_VDD_c_121_n N_A_c_389_n 4.41003e-19
cc_140 N_VDD_c_135_p N_A_c_389_n 6.39485e-19
cc_141 N_SELI_c_189_n N_SEL_c_253_n 8.93041e-19
cc_142 N_SELI_c_192_n N_SEL_c_253_n 3.46631e-19
cc_143 N_SELI_c_209_n N_SEL_c_257_n 0.00339809f
cc_144 N_SELI_c_193_n N_SEL_c_258_n 0.00240446f
cc_145 N_SELI_c_189_n N_SEL_c_259_n 0.0021504f
cc_146 N_SELI_c_192_n N_SEL_c_259_n 0.00339809f
cc_147 N_SELI_c_189_n N_SEL_c_260_n 9.71051e-19
cc_148 N_SELI_c_192_n N_SEL_c_260_n 6.41327e-19
cc_149 N_SELI_c_209_n N_SEL_c_275_n 7.09664e-19
cc_150 N_SELI_c_211_n N_SEL_c_275_n 0.00496695f
cc_151 N_SELI_c_196_n N_SEL_c_275_n 8.74049e-19
cc_152 N_SELI_c_193_n N_SEL_c_262_n 4.99367e-19
cc_153 N_SELI_c_211_n N_SEL_c_262_n 8.86313e-19
cc_154 N_SELI_c_196_n N_SEL_c_262_n 0.00491002f
cc_155 N_SELI_c_193_n N_SEL_c_263_n 0.00165721f
cc_156 N_SELI_c_209_n N_SEL_c_263_n 4.70859e-19
cc_157 N_SELI_c_198_n N_SEL_c_263_n 9.36901e-19
cc_158 N_SELI_c_231_p N_SEL_c_263_n 7.85443e-19
cc_159 N_SELI_c_189_n N_SEL_c_265_n 2.46723e-19
cc_160 N_SELI_c_209_n N_SEL_c_265_n 2.46502e-19
cc_161 N_SELI_c_199_n N_SEL_c_265_n 0.00142585f
cc_162 N_SELI_c_209_n N_SEL_c_266_n 0.00166116f
cc_163 N_SELI_c_198_n N_SEL_c_266_n 7.57935e-19
cc_164 N_SELI_XI5.X0_CG N_B_XI5.X0_PGS 4.34645e-19
cc_165 N_SELI_c_211_n N_B_XI5.X0_PGS 6.90642e-19
cc_166 N_SELI_c_189_n N_B_XI3.X0_PGS 2.37944e-19
cc_167 N_SELI_c_192_n N_B_XI3.X0_PGS 3.60699e-19
cc_168 N_SELI_c_211_n N_B_XI3.X0_PGS 5.45575e-19
cc_169 N_SELI_c_192_n N_B_c_326_n 3.87281e-19
cc_170 N_SELI_c_192_n N_B_c_336_n 5.40503e-19
cc_171 N_SELI_c_192_n B 0.0012892f
cc_172 N_SELI_c_192_n N_B_c_328_n 0.00106294f
cc_173 N_SELI_c_189_n N_Z_c_352_n 5.41397e-19
cc_174 N_SELI_c_193_n N_Z_c_352_n 0.00205681f
cc_175 N_SELI_c_209_n N_Z_c_352_n 0.00246976f
cc_176 N_SELI_c_211_n N_Z_c_352_n 9.16045e-19
cc_177 N_SELI_c_188_n N_A_XI4.X0_PGS 4.5346e-19
cc_178 N_SELI_c_196_n N_A_XI4.X0_PGS 0.00276355f
cc_179 N_SELI_c_196_n N_A_c_389_n 2.00604e-19
cc_180 N_SEL_c_254_n N_B_XI3.X0_PGS 2.04953e-19
cc_181 N_SEL_c_305_p N_B_XI3.X0_PGS 4.64062e-19
cc_182 N_SEL_c_257_n N_B_XI3.X0_PGS 8.04174e-19
cc_183 N_SEL_c_260_n N_B_XI3.X0_PGS 0.00100354f
cc_184 N_SEL_c_275_n N_B_XI3.X0_PGS 0.00142122f
cc_185 N_SEL_c_257_n N_B_c_344_n 2.97958e-19
cc_186 N_SEL_c_260_n N_B_c_344_n 3.50453e-19
cc_187 N_SEL_c_260_n N_B_c_328_n 9.99041e-19
cc_188 N_SEL_c_258_n N_Z_c_352_n 0.00187327f
cc_189 N_SEL_c_274_n N_Z_c_352_n 0.00194252f
cc_190 N_SEL_c_275_n N_Z_c_352_n 9.12105e-19
cc_191 N_SEL_c_262_n N_Z_c_352_n 9.02042e-19
cc_192 N_SEL_c_263_n N_Z_c_352_n 8.60225e-19
cc_193 N_SEL_c_265_n N_Z_c_352_n 0.0021646f
cc_194 N_SEL_c_266_n N_Z_c_352_n 8.38981e-19
cc_195 N_SEL_XI4.X0_CG N_A_XI4.X0_PGS 4.42555e-19
cc_196 N_SEL_c_262_n N_A_XI4.X0_PGS 0.00276355f
cc_197 N_SEL_c_258_n A 7.0885e-19
cc_198 N_SEL_c_262_n A 4.56568e-19
cc_199 N_SEL_XI4.X0_CG N_A_c_389_n 0.00234241f
cc_200 N_SEL_c_258_n N_A_c_389_n 4.99367e-19
cc_201 N_SEL_c_262_n N_A_c_389_n 0.0014909f
cc_202 N_B_XI5.X0_PGS N_A_XI4.X0_PGS 0.00137535f
*
.ends
*
*
.subckt MUXI2_HPNW4 A B S0 Y VDD VSS
xgate (VSS VDD S0 B Y A) G3_MUXI2_N1
.ends
*
* File: G2_NAND2_N1.pex.netlist
* Created: Tue Feb 22 16:31:07 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NAND2_N1_VSS 2 4 6 8 10 20 23 45 50 59 68 69 70 Vss
c27 70 Vss 7.84263e-19
c28 69 Vss 0.00114439f
c29 59 Vss 0.00441797f
c30 50 Vss 5.92201e-19
c31 45 Vss 0.00559837f
c32 38 Vss 0.0299355f
c33 37 Vss 0.0299355f
c34 32 Vss 0.105919f
c35 27 Vss 0.0688517f
c36 23 Vss 6.52493e-20
c37 21 Vss 0.0348456f
c38 20 Vss 0.064644f
c39 10 Vss 0.0834601f
c40 8 Vss 0.0831275f
c41 6 Vss 0.0830428f
c42 4 Vss 0.0828837f
c43 2 Vss 0.00278021f
r44 69 71 0.652036
r45 69 70 1.66714
r46 63 70 0.652036
r47 63 68 9.12761
r48 50 59 1.16709
r49 50 71 2.16729
r50 45 68 4.87639
r51 33 38 0.494161
r52 32 34 0.652036
r53 32 33 2.9175
r54 29 38 0.128424
r55 28 37 0.494161
r56 27 38 0.494161
r57 27 28 2.8008
r58 24 37 0.128424
r59 23 59 0.238214
r60 21 23 1.4004
r61 20 37 0.494161
r62 20 23 1.5171
r63 17 21 0.652036
r64 10 34 2.5674
r65 8 29 2.5674
r66 6 17 2.5674
r67 4 24 2.5674
r68 2 45 1.16709
.ends

.subckt PM_G2_NAND2_N1_VDD 2 4 6 15 17 31 33 34 35 42 44 50 Vss
c43 50 Vss 0.00511687f
c44 42 Vss 0.00686567f
c45 40 Vss 0.00174586f
c46 35 Vss 0.00426091f
c47 34 Vss 8.36616e-19
c48 33 Vss 0.00735566f
c49 31 Vss 0.00189708f
c50 17 Vss 0.184529f
c51 15 Vss 0.0364084f
c52 6 Vss 0.00252742f
c53 4 Vss 0.00226556f
c54 2 Vss 0.0989662f
r55 40 44 0.326018
r56 40 42 4.83471
r57 39 42 7.002
r58 37 50 1.16709
r59 35 39 0.655813
r60 35 37 2.04225
r61 33 44 0.326018
r62 33 34 10.3363
r63 29 34 0.652036
r64 29 31 4.83471
r65 17 50 0.50025
r66 15 17 5.11257
r67 12 15 0.652541
r68 6 42 1.16709
r69 4 31 1.16709
r70 2 12 3.2676
.ends

.subckt PM_G2_NAND2_N1_A 2 4 13 18 21 26 31 Vss
c21 31 Vss 0.00366686f
c22 26 Vss 0.00318863f
c23 18 Vss 0.00132825f
c24 13 Vss 0.0578401f
c25 2 Vss 0.0573541f
r26 23 31 1.16709
r27 21 23 1.91721
r28 18 26 1.16709
r29 18 21 2.9175
r30 13 31 0.50025
r31 10 26 0.50025
r32 4 13 1.80885
r33 2 10 1.80885
.ends

.subckt PM_G2_NAND2_N1_Z 2 4 25 28 Vss
c25 25 Vss 0.00107312f
c26 4 Vss 0.00148239f
c27 2 Vss 0.00149062f
r28 28 30 4.58464
r29 25 28 4.58464
r30 4 30 1.16709
r31 2 25 1.16709
.ends

.subckt PM_G2_NAND2_N1_B 2 4 10 11 14 18 21 Vss
c24 18 Vss 1.08854e-19
c25 14 Vss 0.147604f
c26 11 Vss 0.0356774f
c27 10 Vss 0.286243f
c28 2 Vss 0.174968f
r29 18 21 0.0416786
r30 14 18 1.16709
r31 12 14 2.8008
r32 10 12 0.652036
r33 10 11 8.92755
r34 7 11 0.652036
r35 4 14 3.0342
r36 2 7 5.835
.ends

.subckt G2_NAND2_N1  VSS VDD A Z B
*
* B	B
* Z	Z
* A	A
* VDD	VDD
* VSS	VSS
XI7.X0 N_Z_XI7.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_B_XI7.X0_PGS N_VSS_XI7.X0_S
+ TIGFET_HPNW4
XI8.X0 N_Z_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGS
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI9.X0 N_Z_XI8.X0_D N_VSS_XI9.X0_PGD N_B_XI9.X0_CG N_VSS_XI9.X0_PGS
+ N_VDD_XI9.X0_S TIGFET_HPNW4
*
x_PM_G2_NAND2_N1_VSS N_VSS_XI7.X0_S N_VSS_XI8.X0_PGD N_VSS_XI8.X0_PGS
+ N_VSS_XI9.X0_PGD N_VSS_XI9.X0_PGS N_VSS_c_6_p N_VSS_c_18_p N_VSS_c_1_p
+ N_VSS_c_4_p N_VSS_c_5_p VSS N_VSS_c_9_p N_VSS_c_10_p Vss PM_G2_NAND2_N1_VSS
x_PM_G2_NAND2_N1_VDD N_VDD_XI7.X0_PGD N_VDD_XI8.X0_S N_VDD_XI9.X0_S N_VDD_c_61_p
+ N_VDD_c_54_p N_VDD_c_29_n N_VDD_c_33_n N_VDD_c_37_n N_VDD_c_57_p N_VDD_c_38_n
+ VDD N_VDD_c_43_p Vss PM_G2_NAND2_N1_VDD
x_PM_G2_NAND2_N1_A N_A_XI7.X0_CG N_A_XI8.X0_CG N_A_c_71_n N_A_c_72_n A
+ N_A_c_79_n N_A_c_75_n Vss PM_G2_NAND2_N1_A
x_PM_G2_NAND2_N1_Z N_Z_XI7.X0_D N_Z_XI8.X0_D N_Z_c_94_n Z Vss PM_G2_NAND2_N1_Z
x_PM_G2_NAND2_N1_B N_B_XI7.X0_PGS N_B_XI9.X0_CG N_B_c_117_n N_B_c_119_n
+ N_B_c_123_n N_B_c_127_n B Vss PM_G2_NAND2_N1_B
cc_1 N_VSS_c_1_p N_VDD_XI8.X0_S 0.00136022f
cc_2 N_VSS_XI8.X0_PGS N_VDD_c_29_n 4.05134e-19
cc_3 N_VSS_c_1_p N_VDD_c_29_n 0.00385472f
cc_4 N_VSS_c_4_p N_VDD_c_29_n 0.00232594f
cc_5 N_VSS_c_5_p N_VDD_c_29_n 0.00101015f
cc_6 N_VSS_c_6_p N_VDD_c_33_n 0.00171596f
cc_7 N_VSS_c_4_p N_VDD_c_33_n 0.00161703f
cc_8 N_VSS_c_5_p N_VDD_c_33_n 2.03837e-19
cc_9 N_VSS_c_9_p N_VDD_c_33_n 0.00286543f
cc_10 N_VSS_c_10_p N_VDD_c_37_n 0.00103397f
cc_11 N_VSS_XI9.X0_PGS N_VDD_c_38_n 4.47716e-19
cc_12 N_VSS_c_1_p N_VDD_c_38_n 2.23518e-19
cc_13 N_VSS_c_4_p N_VDD_c_38_n 5.24284e-19
cc_14 N_VSS_c_5_p N_A_c_71_n 0.00234241f
cc_15 N_VSS_c_1_p N_A_c_72_n 0.00297841f
cc_16 N_VSS_c_4_p N_A_c_72_n 8.12473e-19
cc_17 N_VSS_c_5_p N_A_c_72_n 5.42695e-19
cc_18 N_VSS_c_18_p N_A_c_75_n 7.84334e-19
cc_19 N_VSS_c_4_p N_A_c_75_n 4.56568e-19
cc_20 N_VSS_c_5_p N_A_c_75_n 0.00184767f
cc_21 N_VSS_XI7.X0_S N_Z_XI7.X0_D 3.43419e-19
cc_22 N_VSS_c_1_p N_Z_XI7.X0_D 3.48267e-19
cc_23 N_VSS_XI7.X0_S N_Z_c_94_n 3.48267e-19
cc_24 N_VSS_c_1_p N_Z_c_94_n 0.00178967f
cc_25 N_VSS_XI8.X0_PGD N_B_c_117_n 6.72196e-19
cc_26 N_VSS_XI9.X0_PGD N_B_c_117_n 6.72196e-19
cc_27 N_VSS_XI8.X0_PGS N_B_c_119_n 7.91098e-19
cc_28 N_VDD_XI7.X0_PGD N_A_XI7.X0_CG 4.91184e-19
cc_29 N_VDD_XI7.X0_PGD N_A_c_79_n 2.88617e-19
cc_30 N_VDD_c_43_p N_A_c_79_n 7.96439e-19
cc_31 N_VDD_c_33_n N_A_c_75_n 2.29043e-19
cc_32 N_VDD_c_43_p N_Z_XI7.X0_D 0.00132057f
cc_33 N_VDD_XI8.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_34 N_VDD_XI9.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_35 N_VDD_c_29_n N_Z_XI8.X0_D 3.48267e-19
cc_36 N_VDD_c_33_n N_Z_XI8.X0_D 3.7884e-19
cc_37 N_VDD_c_38_n N_Z_XI8.X0_D 3.48267e-19
cc_38 N_VDD_XI7.X0_PGD N_Z_c_94_n 3.00781e-19
cc_39 N_VDD_XI8.X0_S N_Z_c_94_n 3.48267e-19
cc_40 N_VDD_XI9.X0_S N_Z_c_94_n 3.48267e-19
cc_41 N_VDD_c_54_p N_Z_c_94_n 7.07078e-19
cc_42 N_VDD_c_29_n N_Z_c_94_n 5.69026e-19
cc_43 N_VDD_c_33_n N_Z_c_94_n 7.07375e-19
cc_44 N_VDD_c_57_p N_Z_c_94_n 0.00174191f
cc_45 N_VDD_c_38_n N_Z_c_94_n 0.00291831f
cc_46 N_VDD_c_43_p N_Z_c_94_n 8.835e-19
cc_47 N_VDD_XI7.X0_PGD N_B_XI7.X0_PGS 0.00320747f
cc_48 N_VDD_c_61_p N_B_c_117_n 0.0097987f
cc_49 N_VDD_c_38_n N_B_c_117_n 2.48119e-19
cc_50 N_VDD_c_33_n N_B_c_123_n 4.73957e-19
cc_51 N_VDD_c_57_p N_B_c_123_n 3.81676e-19
cc_52 N_VDD_c_38_n N_B_c_123_n 0.001001f
cc_53 N_VDD_c_43_p N_B_c_123_n 0.00150149f
cc_54 N_VDD_c_33_n N_B_c_127_n 4.10393e-19
cc_55 N_VDD_c_57_p N_B_c_127_n 5.19718e-19
cc_56 N_VDD_c_38_n N_B_c_127_n 0.00144738f
cc_57 N_VDD_c_43_p N_B_c_127_n 3.81676e-19
cc_58 N_A_c_72_n N_Z_c_94_n 0.00754545f
cc_59 N_A_c_79_n N_Z_c_94_n 9.58524e-19
cc_60 N_A_c_75_n N_Z_c_94_n 9.18163e-19
cc_61 N_A_XI7.X0_CG N_B_XI7.X0_PGS 4.5346e-19
cc_62 N_A_c_72_n N_B_XI7.X0_PGS 2.82086e-19
cc_63 N_A_c_79_n N_B_XI7.X0_PGS 5.70584e-19
cc_64 N_A_c_72_n N_B_c_117_n 3.21972e-19
cc_65 N_A_c_79_n N_B_c_117_n 0.0014179f
cc_66 N_A_c_75_n N_B_c_117_n 0.00112482f
cc_67 N_A_c_75_n N_B_c_123_n 9.27569e-19
cc_68 N_Z_c_94_n N_B_c_117_n 3.90525e-19
cc_69 N_Z_c_94_n N_B_c_123_n 9.49424e-19
cc_70 N_Z_c_94_n N_B_c_127_n 0.00147334f
*
.ends
*
*
.subckt NAND2_HPNW4 A B Y VDD VSS
xgate (VSS VDD A Y B) G2_NAND2_N1
.ends
*
* File: G2_NOR2_N1.pex.netlist
* Created: Mon Feb 28 09:28:35 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NOR2_N1_VSS 2 4 6 16 18 31 36 41 50 61 62 66 67 72 79 80 Vss
c43 80 Vss 3.75522e-19
c44 79 Vss 0.00223955f
c45 74 Vss 0.00269784f
c46 72 Vss 0.00694708f
c47 67 Vss 8.20725e-19
c48 66 Vss 0.00177669f
c49 62 Vss 6.45375e-19
c50 61 Vss 0.00385292f
c51 50 Vss 0.00491203f
c52 41 Vss 7.10513e-22
c53 36 Vss 9.27479e-19
c54 31 Vss 0.00114656f
c55 18 Vss 0.0881492f
c56 16 Vss 6.95992e-20
c57 6 Vss 0.00202759f
c58 4 Vss 0.0834348f
c59 2 Vss 0.00226843f
r60 78 79 4.16786
r61 74 78 0.655813
r62 73 80 0.494161
r63 72 79 0.652036
r64 72 73 10.1279
r65 68 80 0.128424
r66 66 80 0.494161
r67 66 67 4.37625
r68 59 67 0.652036
r69 59 61 8.46075
r70 58 62 0.655813
r71 58 61 4.87639
r72 41 74 1.82344
r73 36 50 1.16709
r74 36 68 2.16729
r75 31 62 1.82344
r76 16 50 0.238214
r77 16 18 2.04225
r78 12 18 0.0685365
r79 6 41 1.16709
r80 4 12 2.5674
r81 2 31 1.16709
.ends

.subckt PM_G2_NOR2_N1_VDD 2 4 6 8 10 27 29 45 47 48 52 54 55 57 60 64 66 72 78
+ Vss
c51 78 Vss 0.0058262f
c52 72 Vss 0.00492692f
c53 66 Vss 3.56526e-19
c54 64 Vss 9.96234e-19
c55 60 Vss 0.00134431f
c56 55 Vss 8.63545e-19
c57 54 Vss 0.0060792f
c58 52 Vss 0.0016605f
c59 49 Vss 0.00173366f
c60 48 Vss 0.00489508f
c61 47 Vss 0.00194735f
c62 45 Vss 0.00746951f
c63 37 Vss 0.127438f
c64 29 Vss 7.35265e-20
c65 27 Vss 0.0346129f
c66 26 Vss 0.101192f
c67 10 Vss 0.0842957f
c68 8 Vss 0.0823812f
c69 6 Vss 0.00220559f
c70 4 Vss 0.0830779f
c71 2 Vss 0.0842392f
r72 72 75 0.05
r73 64 78 1.16709
r74 62 64 2.16729
r75 60 75 1.16709
r76 58 60 2.20896
r77 55 57 9.04425
r78 54 62 0.652036
r79 54 57 1.12532
r80 50 66 0.0828784
r81 50 52 1.82344
r82 48 58 0.652036
r83 48 49 4.37625
r84 47 55 0.652036
r85 46 66 0.551426
r86 46 47 4.16786
r87 45 66 0.551426
r88 44 49 0.652036
r89 44 45 13.3371
r90 36 72 0.262036
r91 36 37 2.26917
r92 33 36 2.26917
r93 29 78 0.238214
r94 27 29 1.5171
r95 26 30 0.652036
r96 26 29 1.4004
r97 23 27 0.652036
r98 20 37 0.00605528
r99 17 33 0.00605528
r100 10 30 2.5674
r101 8 23 2.5674
r102 6 52 1.16709
r103 4 17 2.5674
r104 2 20 2.5674
.ends

.subckt PM_G2_NOR2_N1_B 2 4 10 13 18 21 26 31 Vss
c25 31 Vss 0.00183593f
c26 26 Vss 0.00362926f
c27 18 Vss 9.68961e-19
c28 13 Vss 0.057478f
c29 10 Vss 6.74849e-20
c30 2 Vss 0.0576626f
r31 23 31 1.16709
r32 21 23 2.20896
r33 18 26 1.16709
r34 18 21 2.62575
r35 13 31 0.50025
r36 10 26 0.50025
r37 4 13 1.80885
r38 2 10 1.80885
.ends

.subckt PM_G2_NOR2_N1_Z 2 4 25 28 Vss
c21 25 Vss 0.00301088f
c22 4 Vss 0.00148239f
c23 2 Vss 0.0021264f
r24 28 30 3.12589
r25 25 28 6.04339
r26 4 30 1.16709
r27 2 25 1.16709
.ends

.subckt PM_G2_NOR2_N1_A 2 4 10 11 14 20 Vss
c18 20 Vss 2.48297e-19
c19 14 Vss 0.116468f
c20 11 Vss 0.0348164f
c21 10 Vss 0.273262f
c22 2 Vss 0.14291f
r23 20 26 1.16709
r24 14 26 0.05
r25 12 14 1.6338
r26 10 12 0.652036
r27 10 11 8.92755
r28 7 11 0.652036
r29 4 14 3.0342
r30 2 7 4.668
.ends

.subckt G2_NOR2_N1  VSS VDD B Z A
*
* A	A
* Z	Z
* B	B
* VDD	VDD
* VSS	VSS
XI2.X0 N_Z_XI2.X0_D N_VDD_XI2.X0_PGD N_B_XI2.X0_CG N_VDD_XI2.X0_PGS
+ N_VSS_XI2.X0_S TIGFET_HPNW4
XI0.X0 N_Z_XI0.X0_D N_VSS_XI0.X0_PGD N_B_XI0.X0_CG N_A_XI0.X0_PGS N_VDD_XI0.X0_S
+ TIGFET_HPNW4
XI1.X0 N_Z_XI0.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
*
x_PM_G2_NOR2_N1_VSS N_VSS_XI2.X0_S N_VSS_XI0.X0_PGD N_VSS_XI1.X0_S N_VSS_c_31_p
+ N_VSS_c_2_p N_VSS_c_4_p N_VSS_c_7_p N_VSS_c_37_p N_VSS_c_8_p VSS N_VSS_c_6_p
+ N_VSS_c_16_p N_VSS_c_19_p N_VSS_c_17_p N_VSS_c_22_p N_VSS_c_18_p Vss
+ PM_G2_NOR2_N1_VSS
x_PM_G2_NOR2_N1_VDD N_VDD_XI2.X0_PGD N_VDD_XI2.X0_PGS N_VDD_XI0.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_c_45_n N_VDD_c_90_p N_VDD_c_46_n
+ N_VDD_c_50_n N_VDD_c_53_n N_VDD_c_55_n N_VDD_c_56_n N_VDD_c_62_n VDD
+ N_VDD_c_72_p N_VDD_c_63_n N_VDD_c_66_n N_VDD_c_69_p N_VDD_c_67_n Vss
+ PM_G2_NOR2_N1_VDD
x_PM_G2_NOR2_N1_B N_B_XI2.X0_CG N_B_XI0.X0_CG N_B_c_104_n N_B_c_95_n N_B_c_96_n
+ B N_B_c_99_n N_B_c_100_n Vss PM_G2_NOR2_N1_B
x_PM_G2_NOR2_N1_Z N_Z_XI2.X0_D N_Z_XI0.X0_D N_Z_c_124_n Z Vss PM_G2_NOR2_N1_Z
x_PM_G2_NOR2_N1_A N_A_XI0.X0_PGS N_A_XI1.X0_CG N_A_c_141_n N_A_c_145_n
+ N_A_c_147_n A Vss PM_G2_NOR2_N1_A
cc_1 N_VSS_XI0.X0_PGD N_VDD_XI1.X0_PGD 0.00180308f
cc_2 N_VSS_c_2_p N_VDD_c_45_n 0.00180308f
cc_3 N_VSS_XI2.X0_S N_VDD_c_46_n 9.5668e-19
cc_4 N_VSS_c_4_p N_VDD_c_46_n 0.00165395f
cc_5 VSS N_VDD_c_46_n 0.00476397f
cc_6 N_VSS_c_6_p N_VDD_c_46_n 0.00186257f
cc_7 N_VSS_c_7_p N_VDD_c_50_n 4.43871e-19
cc_8 N_VSS_c_8_p N_VDD_c_50_n 3.66936e-19
cc_9 VSS N_VDD_c_50_n 0.00285866f
cc_10 N_VSS_XI2.X0_S N_VDD_c_53_n 3.7884e-19
cc_11 N_VSS_c_4_p N_VDD_c_53_n 0.00104703f
cc_12 N_VSS_c_4_p N_VDD_c_55_n 7.47067e-19
cc_13 N_VSS_c_2_p N_VDD_c_56_n 3.37151e-19
cc_14 N_VSS_c_7_p N_VDD_c_56_n 0.00141228f
cc_15 N_VSS_c_8_p N_VDD_c_56_n 0.00112249f
cc_16 N_VSS_c_16_p N_VDD_c_56_n 0.0034844f
cc_17 N_VSS_c_17_p N_VDD_c_56_n 0.00588723f
cc_18 N_VSS_c_18_p N_VDD_c_56_n 7.74609e-19
cc_19 N_VSS_c_19_p N_VDD_c_62_n 0.00106075f
cc_20 N_VSS_c_7_p N_VDD_c_63_n 0.00106112f
cc_21 N_VSS_c_8_p N_VDD_c_63_n 3.95933e-19
cc_22 N_VSS_c_22_p N_VDD_c_63_n 3.86251e-19
cc_23 VSS N_VDD_c_66_n 0.00116512f
cc_24 N_VSS_c_7_p N_VDD_c_67_n 3.44698e-19
cc_25 N_VSS_c_8_p N_VDD_c_67_n 7.95135e-19
cc_26 N_VSS_c_8_p N_B_c_95_n 0.00234321f
cc_27 N_VSS_c_7_p N_B_c_96_n 8.39582e-19
cc_28 N_VSS_c_8_p N_B_c_96_n 5.42695e-19
cc_29 VSS N_B_c_96_n 0.00148607f
cc_30 N_VSS_c_8_p N_B_c_99_n 2.00604e-19
cc_31 N_VSS_c_31_p N_B_c_100_n 8.37306e-19
cc_32 N_VSS_c_7_p N_B_c_100_n 4.56568e-19
cc_33 N_VSS_c_8_p N_B_c_100_n 0.00173573f
cc_34 N_VSS_XI2.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_35 N_VSS_c_4_p N_Z_XI2.X0_D 3.48267e-19
cc_36 N_VSS_XI1.X0_S N_Z_XI0.X0_D 3.43419e-19
cc_37 N_VSS_c_37_p N_Z_XI0.X0_D 3.48267e-19
cc_38 N_VSS_c_4_p N_Z_c_124_n 8.89782e-19
cc_39 N_VSS_c_37_p N_Z_c_124_n 6.0686e-19
cc_40 VSS N_Z_c_124_n 4.63431e-19
cc_41 N_VSS_c_17_p N_Z_c_124_n 2.55365e-19
cc_42 N_VSS_XI0.X0_PGD N_A_c_141_n 9.39677e-19
cc_43 N_VSS_c_2_p N_A_c_141_n 2.16729e-19
cc_44 N_VDD_c_69_p N_B_XI2.X0_CG 0.00237871f
cc_45 N_VDD_c_69_p N_B_c_104_n 0.0010681f
cc_46 N_VDD_c_46_n N_B_c_96_n 0.0025037f
cc_47 N_VDD_c_72_p N_B_c_96_n 7.41679e-19
cc_48 N_VDD_c_69_p N_B_c_96_n 5.48133e-19
cc_49 N_VDD_c_46_n N_B_c_99_n 4.9897e-19
cc_50 N_VDD_c_72_p N_B_c_99_n 4.91501e-19
cc_51 N_VDD_c_69_p N_B_c_99_n 0.00150793f
cc_52 N_VDD_c_46_n N_B_c_100_n 3.66936e-19
cc_53 N_VDD_c_69_p N_B_c_100_n 2.00604e-19
cc_54 N_VDD_XI0.X0_S N_Z_XI0.X0_D 3.43419e-19
cc_55 N_VDD_c_55_n N_Z_XI0.X0_D 3.72199e-19
cc_56 N_VDD_c_56_n N_Z_XI0.X0_D 3.7884e-19
cc_57 N_VDD_XI0.X0_S N_Z_c_124_n 3.48267e-19
cc_58 N_VDD_c_46_n N_Z_c_124_n 5.1034e-19
cc_59 N_VDD_c_55_n N_Z_c_124_n 7.89245e-19
cc_60 N_VDD_c_56_n N_Z_c_124_n 5.36364e-19
cc_61 N_VDD_XI2.X0_PGD N_A_c_141_n 5.10213e-19
cc_62 N_VDD_XI1.X0_PGD N_A_c_141_n 2.48727e-19
cc_63 N_VDD_XI2.X0_PGS N_A_c_145_n 6.4837e-19
cc_64 N_VDD_c_46_n N_A_c_145_n 3.16598e-19
cc_65 N_VDD_c_90_p N_A_c_147_n 8.9931e-19
cc_66 N_VDD_c_63_n N_A_c_147_n 4.91217e-19
cc_67 N_VDD_c_67_n N_A_c_147_n 0.00320668f
cc_68 N_VDD_c_63_n A 6.1931e-19
cc_69 N_VDD_c_67_n A 4.56568e-19
cc_70 N_B_c_96_n N_Z_c_124_n 0.00744925f
cc_71 N_B_c_99_n N_Z_c_124_n 9.58524e-19
cc_72 N_B_c_100_n N_Z_c_124_n 8.92526e-19
cc_73 N_B_c_95_n N_A_XI0.X0_PGS 4.5346e-19
cc_74 N_B_c_100_n N_A_XI0.X0_PGS 7.86826e-19
cc_75 N_B_c_99_n N_A_c_141_n 9.25308e-19
cc_76 N_B_c_100_n N_A_c_147_n 7.50183e-19
cc_77 N_Z_c_124_n N_A_c_141_n 9.72643e-19
cc_78 N_Z_c_124_n N_A_c_147_n 9.67259e-19
cc_79 N_Z_c_124_n A 0.00155484f
*
.ends
*
*
.subckt NOR2_HPNW4 A B Y VDD VSS
xgate (VSS VDD B Y A) G2_NOR2_N1
.ends
*
* File: G2_OAI21_N1.pex.netlist
* Created: Wed Feb 23 15:42:41 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_OAI21_N1_VSS 2 4 6 8 10 22 29 45 50 55 64 73 74 78 84 86 91 94 Vss
c49 92 Vss 5.73928e-19
c50 91 Vss 0.00675279f
c51 86 Vss 0.00175471f
c52 84 Vss 0.00280649f
c53 79 Vss 0.00136179f
c54 78 Vss 0.00706512f
c55 74 Vss 6.45375e-19
c56 73 Vss 0.00483551f
c57 64 Vss 0.00536833f
c58 55 Vss 1.70165e-19
c59 50 Vss 0.00185649f
c60 45 Vss 0.0012795f
c61 33 Vss 0.0307391f
c62 29 Vss 7.39492e-20
c63 26 Vss 0.101218f
c64 22 Vss 0.0345446f
c65 21 Vss 0.0712517f
c66 10 Vss 0.0820743f
c67 8 Vss 0.0810902f
c68 6 Vss 0.00226958f
c69 4 Vss 0.0806996f
c70 2 Vss 0.00266945f
r71 91 94 0.326018
r72 90 91 13.3371
r73 86 90 0.655813
r74 85 92 0.494161
r75 84 94 0.326018
r76 84 85 4.33457
r77 80 92 0.128424
r78 78 92 0.494161
r79 78 79 10.1696
r80 73 79 0.652036
r81 72 74 0.655813
r82 72 73 13.3371
r83 55 86 1.82344
r84 50 64 1.16709
r85 50 80 2.16729
r86 45 74 1.82344
r87 29 64 0.238214
r88 27 33 0.494161
r89 27 29 1.5171
r90 26 30 0.652036
r91 26 29 1.4004
r92 23 33 0.128424
r93 21 33 0.494161
r94 21 22 2.8008
r95 18 22 0.652036
r96 10 30 2.5674
r97 8 23 2.5674
r98 6 55 1.16709
r99 4 18 2.5674
r100 2 45 1.16709
.ends

.subckt PM_G2_OAI21_N1_VDD 2 4 6 8 38 39 41 43 47 49 51 56 59 65 Vss
c51 65 Vss 0.00591189f
c52 57 Vss 5.34798e-19
c53 56 Vss 0.00857327f
c54 51 Vss 0.00150304f
c55 49 Vss 0.00549985f
c56 47 Vss 0.00136862f
c57 43 Vss 0.00161014f
c58 41 Vss 7.26487e-19
c59 40 Vss 0.00177073f
c60 39 Vss 0.00917963f
c61 38 Vss 0.00784728f
c62 25 Vss 0.085695f
c63 19 Vss 0.0340946f
c64 18 Vss 0.0688517f
c65 8 Vss 0.00226556f
c66 6 Vss 0.0830486f
c67 4 Vss 0.00236553f
c68 2 Vss 0.0834535f
r69 56 59 0.349767
r70 55 56 13.3371
r71 51 59 0.306046
r72 51 53 1.82344
r73 50 57 0.494161
r74 49 55 0.652036
r75 49 50 4.37625
r76 47 65 1.16709
r77 45 57 0.128424
r78 45 47 2.16729
r79 41 43 1.82344
r80 39 57 0.494161
r81 39 40 10.1279
r82 38 41 0.655813
r83 37 40 0.652036
r84 37 38 13.3371
r85 25 65 0.238214
r86 23 25 2.04225
r87 20 23 0.0685365
r88 18 23 0.5835
r89 18 19 2.8008
r90 15 19 0.652036
r91 8 53 1.16709
r92 6 20 2.5674
r93 4 43 1.16709
r94 2 15 2.5674
.ends

.subckt PM_G2_OAI21_N1_B 2 4 10 13 18 21 26 31 Vss
c23 31 Vss 0.00366366f
c24 26 Vss 0.00309808f
c25 18 Vss 6.90549e-19
c26 13 Vss 0.0578401f
c27 2 Vss 0.0576308f
r28 23 31 1.16709
r29 21 23 1.95889
r30 18 26 1.16709
r31 18 21 2.87582
r32 13 31 0.50025
r33 10 26 0.50025
r34 4 13 1.80885
r35 2 10 1.80885
.ends

.subckt PM_G2_OAI21_N1_A 2 4 13 18 26 31 36 43 45 Vss
c43 43 Vss 0.0016451f
c44 36 Vss 0.00277103f
c45 31 Vss 0.00697771f
c46 26 Vss 0.00360766f
c47 18 Vss 0.0860562f
c48 13 Vss 6.71834e-20
c49 4 Vss 0.0575023f
c50 2 Vss 0.0840749f
r51 40 45 0.655813
r52 40 43 9.00257
r53 31 43 1.16709
r54 26 36 1.16709
r55 26 45 4.52212
r56 18 31 0.238214
r57 15 18 1.92555
r58 13 36 0.50025
r59 7 15 0.0685365
r60 4 13 1.80885
r61 2 7 2.5674
.ends

.subckt PM_G2_OAI21_N1_Z 2 4 30 33 Vss
c30 30 Vss 0.00127106f
c31 4 Vss 0.00153036f
c32 2 Vss 0.00148239f
r33 33 35 5.62661
r34 30 33 3.54268
r35 4 35 1.16709
r36 2 30 1.16709
.ends

.subckt PM_G2_OAI21_N1_C 2 4 6 13 14 17 24 27 30 Vss
c30 27 Vss 4.95129e-19
c31 24 Vss 0.0812483f
c32 17 Vss 0.147907f
c33 14 Vss 0.0348316f
c34 13 Vss 0.245605f
c35 4 Vss 0.18102f
c36 2 Vss 0.181207f
r37 27 30 0.0833571
r38 23 24 2.04225
r39 20 24 0.0685365
r40 17 27 1.16709
r41 15 23 0.0685365
r42 15 17 2.8008
r43 13 23 0.5835
r44 13 14 8.92755
r45 10 14 0.652036
r46 6 17 3.0342
r47 4 20 5.835
r48 2 10 5.835
.ends

.subckt G2_OAI21_N1  VSS VDD B A Z C
*
* C	C
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI1.X0 N_Z_XI1.X0_D N_VDD_XI1.X0_PGD N_B_XI1.X0_CG N_C_XI1.X0_PGS N_VSS_XI1.X0_S
+ TIGFET_HPNW4
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_A_XI6.X0_PGS N_VDD_XI6.X0_S
+ TIGFET_HPNW4
XI5.X0 N_Z_XI1.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_C_XI5.X0_PGS N_VSS_XI5.X0_S
+ TIGFET_HPNW4
XI7.X0 N_Z_XI6.X0_D N_VSS_XI7.X0_PGD N_C_XI7.X0_CG N_VSS_XI7.X0_PGS
+ N_VDD_XI7.X0_S TIGFET_HPNW4
*
x_PM_G2_OAI21_N1_VSS N_VSS_XI1.X0_S N_VSS_XI6.X0_PGD N_VSS_XI5.X0_S
+ N_VSS_XI7.X0_PGD N_VSS_XI7.X0_PGS N_VSS_c_22_p N_VSS_c_44_p N_VSS_c_1_p
+ N_VSS_c_23_p N_VSS_c_9_p N_VSS_c_24_p N_VSS_c_2_p N_VSS_c_3_p N_VSS_c_7_p
+ N_VSS_c_12_p N_VSS_c_10_p N_VSS_c_16_p VSS Vss PM_G2_OAI21_N1_VSS
x_PM_G2_OAI21_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI6.X0_S N_VDD_XI5.X0_PGD
+ N_VDD_XI7.X0_S N_VDD_c_50_n N_VDD_c_53_n N_VDD_c_54_n N_VDD_c_55_n
+ N_VDD_c_75_p N_VDD_c_57_n N_VDD_c_60_n N_VDD_c_63_n VDD N_VDD_c_72_p Vss
+ PM_G2_OAI21_N1_VDD
x_PM_G2_OAI21_N1_B N_B_XI1.X0_CG N_B_XI6.X0_CG N_B_c_102_n N_B_c_109_p
+ N_B_c_101_n B N_B_c_105_n N_B_c_107_n Vss PM_G2_OAI21_N1_B
x_PM_G2_OAI21_N1_A N_A_XI6.X0_PGS N_A_XI5.X0_CG N_A_c_139_n N_A_c_149_n
+ N_A_c_125_n N_A_c_127_n N_A_c_131_n A N_A_c_137_n Vss PM_G2_OAI21_N1_A
x_PM_G2_OAI21_N1_Z N_Z_XI1.X0_D N_Z_XI6.X0_D N_Z_c_171_n Z Vss PM_G2_OAI21_N1_Z
x_PM_G2_OAI21_N1_C N_C_XI1.X0_PGS N_C_XI5.X0_PGS N_C_XI7.X0_CG N_C_c_197_n
+ N_C_c_219_n N_C_c_199_n N_C_c_202_n N_C_c_203_n C Vss PM_G2_OAI21_N1_C
cc_1 N_VSS_c_1_p N_VDD_c_50_n 0.00187494f
cc_2 N_VSS_c_2_p N_VDD_c_50_n 0.00510452f
cc_3 N_VSS_c_3_p N_VDD_c_50_n 0.00186257f
cc_4 N_VSS_c_1_p N_VDD_c_53_n 0.0010904f
cc_5 N_VSS_c_2_p N_VDD_c_54_n 0.0014876f
cc_6 N_VSS_c_1_p N_VDD_c_55_n 7.48363e-19
cc_7 N_VSS_c_7_p N_VDD_c_55_n 4.59722e-19
cc_8 N_VSS_XI5.X0_S N_VDD_c_57_n 3.7884e-19
cc_9 N_VSS_c_9_p N_VDD_c_57_n 5.11058e-19
cc_10 N_VSS_c_10_p N_VDD_c_57_n 5.35974e-19
cc_11 N_VSS_c_9_p N_VDD_c_60_n 2.14355e-19
cc_12 N_VSS_c_12_p N_VDD_c_60_n 4.59722e-19
cc_13 N_VSS_c_10_p N_VDD_c_60_n 5.34009e-19
cc_14 N_VSS_c_9_p N_VDD_c_63_n 0.00187494f
cc_15 N_VSS_c_10_p N_VDD_c_63_n 0.00186257f
cc_16 N_VSS_c_16_p N_VDD_c_63_n 0.00730042f
cc_17 N_VSS_c_2_p N_B_c_101_n 5.86846e-19
cc_18 N_VSS_XI6.X0_PGD N_A_XI6.X0_PGS 0.00164631f
cc_19 N_VSS_c_7_p N_A_c_125_n 8.83597e-19
cc_20 N_VSS_c_16_p N_A_c_125_n 4.02032e-19
cc_21 N_VSS_XI6.X0_PGD N_A_c_127_n 3.11814e-19
cc_22 N_VSS_c_22_p N_A_c_127_n 0.00322564f
cc_23 N_VSS_c_23_p N_A_c_127_n 3.44698e-19
cc_24 N_VSS_c_24_p N_A_c_127_n 6.61253e-19
cc_25 N_VSS_c_24_p N_A_c_131_n 3.77503e-19
cc_26 N_VSS_c_23_p A 8.59446e-19
cc_27 N_VSS_c_24_p A 3.44698e-19
cc_28 N_VSS_c_2_p A 0.00272781f
cc_29 N_VSS_c_7_p A 0.00211023f
cc_30 N_VSS_c_16_p A 0.00133784f
cc_31 N_VSS_c_2_p N_A_c_137_n 0.00291082f
cc_32 N_VSS_XI1.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_33 N_VSS_XI5.X0_S N_Z_XI1.X0_D 3.43419e-19
cc_34 N_VSS_c_1_p N_Z_XI1.X0_D 3.48267e-19
cc_35 N_VSS_c_9_p N_Z_XI1.X0_D 3.48267e-19
cc_36 N_VSS_XI1.X0_S N_Z_c_171_n 3.48267e-19
cc_37 N_VSS_XI5.X0_S N_Z_c_171_n 3.48267e-19
cc_38 N_VSS_c_1_p N_Z_c_171_n 5.69026e-19
cc_39 N_VSS_c_9_p N_Z_c_171_n 5.69026e-19
cc_40 N_VSS_c_7_p N_Z_c_171_n 4.84633e-19
cc_41 N_VSS_c_16_p N_Z_c_171_n 4.50981e-19
cc_42 N_VSS_XI6.X0_PGD N_C_c_197_n 6.77138e-19
cc_43 N_VSS_XI7.X0_PGD N_C_c_197_n 6.77138e-19
cc_44 N_VSS_c_44_p N_C_c_199_n 8.9608e-19
cc_45 N_VSS_c_23_p N_C_c_199_n 4.56568e-19
cc_46 N_VSS_c_24_p N_C_c_199_n 0.00315719f
cc_47 N_VSS_XI7.X0_PGS N_C_c_202_n 7.91098e-19
cc_48 N_VSS_c_23_p N_C_c_203_n 5.37794e-19
cc_49 N_VSS_c_24_p N_C_c_203_n 4.56568e-19
cc_50 N_VDD_c_53_n N_B_c_102_n 2.44914e-19
cc_51 N_VDD_c_50_n N_B_c_101_n 0.00216638f
cc_52 N_VDD_c_53_n N_B_c_101_n 2.85486e-19
cc_53 N_VDD_c_50_n N_B_c_105_n 3.66936e-19
cc_54 N_VDD_c_53_n N_B_c_105_n 2.29043e-19
cc_55 N_VDD_c_50_n N_B_c_107_n 4.1997e-19
cc_56 N_VDD_c_72_p N_A_XI5.X0_CG 0.00237871f
cc_57 N_VDD_c_72_p N_A_c_139_n 0.00106215f
cc_58 N_VDD_c_53_n N_A_c_125_n 9.72202e-19
cc_59 N_VDD_c_75_p N_A_c_125_n 7.80108e-19
cc_60 N_VDD_c_63_n N_A_c_125_n 6.23587e-19
cc_61 N_VDD_c_72_p N_A_c_125_n 4.87728e-19
cc_62 N_VDD_c_75_p N_A_c_131_n 4.85469e-19
cc_63 N_VDD_c_63_n N_A_c_131_n 3.66936e-19
cc_64 N_VDD_c_72_p N_A_c_131_n 0.0014909f
cc_65 N_VDD_c_50_n N_A_c_137_n 6.23756e-19
cc_66 N_VDD_c_53_n N_A_c_137_n 2.0345e-19
cc_67 N_VDD_c_53_n N_Z_XI1.X0_D 3.7884e-19
cc_68 N_VDD_XI6.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_69 N_VDD_XI7.X0_S N_Z_XI6.X0_D 3.43419e-19
cc_70 N_VDD_c_55_n N_Z_XI6.X0_D 3.72199e-19
cc_71 N_VDD_c_60_n N_Z_XI6.X0_D 3.72199e-19
cc_72 N_VDD_XI6.X0_S N_Z_c_171_n 3.48267e-19
cc_73 N_VDD_XI7.X0_S N_Z_c_171_n 3.48267e-19
cc_74 N_VDD_c_50_n N_Z_c_171_n 3.87755e-19
cc_75 N_VDD_c_53_n N_Z_c_171_n 6.81554e-19
cc_76 N_VDD_c_55_n N_Z_c_171_n 5.6271e-19
cc_77 N_VDD_c_60_n N_Z_c_171_n 7.76033e-19
cc_78 N_VDD_c_63_n N_Z_c_171_n 0.0010014f
cc_79 N_VDD_c_50_n N_C_XI1.X0_PGS 6.09123e-19
cc_80 N_VDD_c_63_n N_C_XI5.X0_PGS 6.28572e-19
cc_81 N_VDD_XI1.X0_PGD N_C_c_197_n 6.72196e-19
cc_82 N_VDD_XI5.X0_PGD N_C_c_197_n 6.76891e-19
cc_83 N_VDD_c_63_n N_C_c_199_n 4.79801e-19
cc_84 N_VDD_c_63_n N_C_c_203_n 3.46645e-19
cc_85 N_B_c_107_n N_A_c_149_n 8.43061e-19
cc_86 N_B_c_109_p N_A_c_127_n 0.00234241f
cc_87 N_B_c_101_n N_A_c_127_n 5.28799e-19
cc_88 N_B_c_107_n N_A_c_127_n 0.00173494f
cc_89 N_B_c_105_n N_A_c_131_n 8.86454e-19
cc_90 N_B_c_101_n A 0.00306515f
cc_91 N_B_c_107_n A 4.56568e-19
cc_92 N_B_c_101_n N_A_c_137_n 6.59436e-19
cc_93 N_B_c_101_n N_Z_c_171_n 0.00673203f
cc_94 N_B_c_105_n N_Z_c_171_n 9.17696e-19
cc_95 N_B_c_107_n N_Z_c_171_n 9.18163e-19
cc_96 N_B_XI1.X0_CG N_C_XI1.X0_PGS 4.42555e-19
cc_97 N_B_c_105_n N_C_XI1.X0_PGS 0.001089f
cc_98 N_B_c_105_n N_C_c_197_n 6.02551e-19
cc_99 N_B_c_107_n N_C_c_197_n 0.00107456f
cc_100 N_B_c_107_n N_C_c_199_n 9.3196e-19
cc_101 N_A_c_125_n N_Z_c_171_n 0.00382179f
cc_102 A N_Z_c_171_n 0.00134325f
cc_103 N_A_XI5.X0_CG N_C_XI5.X0_PGS 4.42555e-19
cc_104 N_A_c_131_n N_C_XI5.X0_PGS 0.001089f
cc_105 N_A_c_131_n N_C_c_197_n 6.59241e-19
cc_106 N_A_XI6.X0_PGS N_C_c_219_n 7.91098e-19
cc_107 N_A_c_125_n N_C_c_199_n 5.38228e-19
cc_108 N_A_c_127_n N_C_c_199_n 2.62413e-19
cc_109 N_A_c_131_n N_C_c_199_n 0.0021499f
cc_110 N_A_c_125_n N_C_c_203_n 8.10255e-19
cc_111 N_Z_c_171_n N_C_c_197_n 4.9701e-19
cc_112 N_Z_c_171_n N_C_c_199_n 9.61365e-19
cc_113 N_Z_c_171_n N_C_c_203_n 0.00143964f
*
.ends
*
*
.subckt OAI21_HPNW4 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 A0 Y B0) G2_OAI21_N1
.ends
*
* File: G3_OR2_N1.pex.netlist
* Created: Tue Mar  1 11:26:38 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_OR2_N1_VSS 2 4 6 10 12 28 29 36 38 52 57 62 67 76 85 90 91 95 96
+ 101 107 113 115 Vss
c75 115 Vss 3.87529e-19
c76 113 Vss 3.75522e-19
c77 107 Vss 0.00356169f
c78 101 Vss 0.00288979f
c79 96 Vss 8.28047e-19
c80 95 Vss 0.00177669f
c81 91 Vss 6.45375e-19
c82 90 Vss 0.00387778f
c83 85 Vss 0.00483971f
c84 76 Vss 0.00487294f
c85 67 Vss 9.52891e-19
c86 62 Vss 6.68032e-19
c87 57 Vss 8.26459e-19
c88 52 Vss 0.00114656f
c89 38 Vss 0.0883089f
c90 36 Vss 6.95992e-20
c91 29 Vss 0.0339709f
c92 28 Vss 0.0988304f
c93 12 Vss 0.0842992f
c94 10 Vss 0.0825208f
c95 6 Vss 0.00148239f
c96 4 Vss 0.0834348f
c97 2 Vss 0.00226843f
r98 108 115 0.494161
r99 107 109 0.652036
r100 107 108 7.46046
r101 103 115 0.128424
r102 102 113 0.494161
r103 101 115 0.494161
r104 101 102 7.46046
r105 97 113 0.128424
r106 95 113 0.494161
r107 95 96 4.37625
r108 90 96 0.652036
r109 89 91 0.655813
r110 89 90 13.3371
r111 67 85 1.16709
r112 67 109 2.16729
r113 62 103 4.83471
r114 57 76 1.16709
r115 57 97 2.16729
r116 52 91 1.82344
r117 36 76 0.238214
r118 36 38 2.04225
r119 31 85 0.238214
r120 29 31 1.45875
r121 28 32 0.652036
r122 28 31 1.45875
r123 25 29 0.652036
r124 22 38 0.0685365
r125 12 32 2.5674
r126 10 25 2.5674
r127 6 62 1.16709
r128 4 22 2.5674
r129 2 52 1.16709
.ends

.subckt PM_G3_OR2_N1_VDD 2 4 6 8 10 12 14 16 37 39 46 49 70 72 73 77 79 83 87 89
+ 93 95 97 102 103 105 106 107 113 119 124 Vss
c84 124 Vss 0.00429743f
c85 119 Vss 0.00559477f
c86 113 Vss 0.00492664f
c87 107 Vss 2.39889e-19
c88 106 Vss 2.39889e-19
c89 103 Vss 3.56526e-19
c90 102 Vss 0.00314642f
c91 97 Vss 0.00307382f
c92 95 Vss 0.00838282f
c93 93 Vss 5.19372e-19
c94 89 Vss 0.00212525f
c95 87 Vss 4.89903e-19
c96 83 Vss 0.00134401f
c97 79 Vss 0.00561519f
c98 77 Vss 0.0016605f
c99 74 Vss 0.00173366f
c100 73 Vss 0.0048947f
c101 72 Vss 0.00279823f
c102 70 Vss 0.00738679f
c103 57 Vss 0.126882f
c104 47 Vss 0.0348458f
c105 46 Vss 0.1003f
c106 39 Vss 7.35265e-20
c107 37 Vss 0.0346129f
c108 36 Vss 0.100535f
c109 16 Vss 0.00262047f
c110 14 Vss 0.0828904f
c111 12 Vss 0.0825208f
c112 10 Vss 0.0828869f
c113 8 Vss 0.0823812f
c114 6 Vss 0.00220666f
c115 4 Vss 0.0830779f
c116 2 Vss 0.0842392f
r117 113 116 0.05
r118 101 102 4.16786
r119 97 101 0.655813
r120 97 99 1.82344
r121 96 107 0.494161
r122 95 102 0.652036
r123 95 96 10.1279
r124 93 124 1.16709
r125 91 107 0.128424
r126 91 93 2.16729
r127 90 106 0.494161
r128 89 107 0.494161
r129 89 90 4.54296
r130 87 119 1.16709
r131 85 106 0.128424
r132 85 87 2.16729
r133 83 116 1.16709
r134 81 83 2.20896
r135 80 105 0.326018
r136 79 106 0.494161
r137 79 80 10.1696
r138 75 103 0.0828784
r139 75 77 1.82344
r140 73 81 0.652036
r141 73 74 4.37625
r142 72 105 0.326018
r143 71 103 0.551426
r144 71 72 4.16786
r145 70 103 0.551426
r146 69 74 0.652036
r147 69 70 13.3371
r148 56 113 0.262036
r149 56 57 2.26917
r150 53 56 2.26917
r151 49 124 0.238214
r152 47 49 1.45875
r153 46 50 0.652036
r154 46 49 1.45875
r155 43 47 0.652036
r156 39 119 0.238214
r157 37 39 1.5171
r158 36 40 0.652036
r159 36 39 1.4004
r160 33 37 0.652036
r161 30 57 0.00605528
r162 27 53 0.00605528
r163 16 99 1.16709
r164 14 43 2.5674
r165 12 50 2.5674
r166 10 40 2.5674
r167 8 33 2.5674
r168 6 77 1.16709
r169 4 27 2.5674
r170 2 30 2.5674
.ends

.subckt PM_G3_OR2_N1_B 2 4 10 13 18 21 26 31 Vss
c25 31 Vss 0.00183593f
c26 26 Vss 0.00362926f
c27 18 Vss 0.00110935f
c28 13 Vss 0.057478f
c29 10 Vss 6.71834e-20
c30 2 Vss 0.0576626f
r31 23 31 1.16709
r32 21 23 2.08393
r33 18 26 1.16709
r34 18 21 2.75079
r35 13 31 0.50025
r36 10 26 0.50025
r37 4 13 1.80885
r38 2 10 1.80885
.ends

.subckt PM_G3_OR2_N1_NET21 2 4 8 10 21 24 45 53 66 70 Vss
c39 70 Vss 0.00761723f
c40 66 Vss 0.00611981f
c41 53 Vss 0.00155023f
c42 45 Vss 0.00245986f
c43 24 Vss 0.225594f
c44 21 Vss 0.0713786f
c45 19 Vss 0.0247918f
c46 10 Vss 0.0847975f
c47 4 Vss 0.00148239f
c48 2 Vss 0.0021264f
r49 70 74 0.652036
r50 53 66 1.16709
r51 53 74 2.9175
r52 48 70 8.04396
r53 48 50 5.66829
r54 45 48 3.501
r55 27 66 0.0476429
r56 25 27 0.326018
r57 25 27 0.1167
r58 24 28 0.652036
r59 24 27 6.7686
r60 21 66 0.357321
r61 19 27 0.326018
r62 19 21 0.40845
r63 10 28 2.5674
r64 8 21 2.15895
r65 4 50 1.16709
r66 2 45 1.16709
.ends

.subckt PM_G3_OR2_N1_A 2 4 10 11 14 18 Vss
c22 18 Vss 2.95942e-19
c23 14 Vss 0.116245f
c24 11 Vss 0.0348164f
c25 10 Vss 0.273261f
c26 2 Vss 0.142908f
r27 21 27 1.16709
r28 18 21 0.0833571
r29 14 27 0.05
r30 12 14 1.6338
r31 10 12 0.652036
r32 10 11 8.92755
r33 7 11 0.652036
r34 4 14 3.0342
r35 2 7 4.668
.ends

.subckt PM_G3_OR2_N1_Z 2 16 19 Vss
c11 2 Vss 0.00148239f
r12 16 19 0.0364688
r13 2 19 1.16709
.ends

.subckt G3_OR2_N1  VSS VDD B A Z
*
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI2.X0 N_NET21_XI2.X0_D N_VDD_XI2.X0_PGD N_B_XI2.X0_CG N_VDD_XI2.X0_PGS
+ N_VSS_XI2.X0_S TIGFET_HPNW4
XI0.X0 N_NET21_XI0.X0_D N_VSS_XI0.X0_PGD N_B_XI0.X0_CG N_A_XI0.X0_PGS
+ N_VDD_XI0.X0_S TIGFET_HPNW4
XI1.X0 N_NET21_XI0.X0_D N_VDD_XI1.X0_PGD N_A_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI3.X0 N_Z_XI3.X0_D N_VDD_XI3.X0_PGD N_NET21_XI3.X0_CG N_VDD_XI3.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI4.X0 N_Z_XI3.X0_D N_VSS_XI4.X0_PGD N_NET21_XI4.X0_CG N_VSS_XI4.X0_PGS
+ N_VDD_XI4.X0_S TIGFET_HPNW4
*
x_PM_G3_OR2_N1_VSS N_VSS_XI2.X0_S N_VSS_XI0.X0_PGD N_VSS_XI1.X0_S
+ N_VSS_XI4.X0_PGD N_VSS_XI4.X0_PGS N_VSS_c_32_p N_VSS_c_4_p N_VSS_c_51_p
+ N_VSS_c_3_p N_VSS_c_6_p N_VSS_c_9_p N_VSS_c_23_p N_VSS_c_30_p N_VSS_c_10_p
+ N_VSS_c_31_p N_VSS_c_7_p N_VSS_c_8_p N_VSS_c_19_p N_VSS_c_12_p N_VSS_c_20_p
+ N_VSS_c_27_p N_VSS_c_21_p VSS Vss PM_G3_OR2_N1_VSS
x_PM_G3_OR2_N1_VDD N_VDD_XI2.X0_PGD N_VDD_XI2.X0_PGS N_VDD_XI0.X0_S
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI3.X0_PGD N_VDD_XI3.X0_PGS
+ N_VDD_XI4.X0_S N_VDD_c_78_n N_VDD_c_149_p N_VDD_c_79_n N_VDD_c_140_p
+ N_VDD_c_80_n N_VDD_c_84_n N_VDD_c_88_n N_VDD_c_90_n N_VDD_c_91_n N_VDD_c_124_p
+ N_VDD_c_97_n N_VDD_c_100_n N_VDD_c_104_n N_VDD_c_107_n N_VDD_c_156_p
+ N_VDD_c_112_n N_VDD_c_114_n VDD N_VDD_c_115_n N_VDD_c_116_n N_VDD_c_121_p
+ N_VDD_c_117_n N_VDD_c_119_n Vss PM_G3_OR2_N1_VDD
x_PM_G3_OR2_N1_B N_B_XI2.X0_CG N_B_XI0.X0_CG N_B_c_169_n N_B_c_160_n N_B_c_161_n
+ B N_B_c_164_n N_B_c_165_n Vss PM_G3_OR2_N1_B
x_PM_G3_OR2_N1_NET21 N_NET21_XI2.X0_D N_NET21_XI0.X0_D N_NET21_XI3.X0_CG
+ N_NET21_XI4.X0_CG N_NET21_c_203_n N_NET21_c_190_n N_NET21_c_191_n
+ N_NET21_c_195_n N_NET21_c_212_n N_NET21_c_197_n Vss PM_G3_OR2_N1_NET21
x_PM_G3_OR2_N1_A N_A_XI0.X0_PGS N_A_XI1.X0_CG N_A_c_224_n N_A_c_228_n
+ N_A_c_230_n A Vss PM_G3_OR2_N1_A
x_PM_G3_OR2_N1_Z N_Z_XI3.X0_D Z N_Z_c_248_n Vss PM_G3_OR2_N1_Z
cc_1 N_VSS_XI0.X0_PGD N_VDD_XI1.X0_PGD 0.00175996f
cc_2 N_VSS_XI4.X0_PGD N_VDD_XI3.X0_PGD 0.00168578f
cc_3 N_VSS_c_3_p N_VDD_c_78_n 0.00175996f
cc_4 N_VSS_c_4_p N_VDD_c_79_n 0.00168578f
cc_5 N_VSS_XI2.X0_S N_VDD_c_80_n 9.5668e-19
cc_6 N_VSS_c_6_p N_VDD_c_80_n 0.00165395f
cc_7 N_VSS_c_7_p N_VDD_c_80_n 0.00519974f
cc_8 N_VSS_c_8_p N_VDD_c_80_n 0.00186257f
cc_9 N_VSS_c_9_p N_VDD_c_84_n 4.43871e-19
cc_10 N_VSS_c_10_p N_VDD_c_84_n 3.66936e-19
cc_11 N_VSS_c_7_p N_VDD_c_84_n 0.00303537f
cc_12 N_VSS_c_12_p N_VDD_c_84_n 0.00106607f
cc_13 N_VSS_XI2.X0_S N_VDD_c_88_n 3.7884e-19
cc_14 N_VSS_c_6_p N_VDD_c_88_n 0.00104703f
cc_15 N_VSS_c_6_p N_VDD_c_90_n 7.47067e-19
cc_16 N_VSS_c_3_p N_VDD_c_91_n 3.37151e-19
cc_17 N_VSS_c_9_p N_VDD_c_91_n 0.00161703f
cc_18 N_VSS_c_10_p N_VDD_c_91_n 2.03837e-19
cc_19 N_VSS_c_19_p N_VDD_c_91_n 0.0034844f
cc_20 N_VSS_c_20_p N_VDD_c_91_n 0.00432568f
cc_21 N_VSS_c_21_p N_VDD_c_91_n 7.74609e-19
cc_22 N_VSS_c_9_p N_VDD_c_97_n 8.45115e-19
cc_23 N_VSS_c_23_p N_VDD_c_97_n 3.93845e-19
cc_24 N_VSS_c_10_p N_VDD_c_97_n 3.95933e-19
cc_25 N_VSS_c_23_p N_VDD_c_100_n 5.01863e-19
cc_26 N_VSS_c_20_p N_VDD_c_100_n 0.00137553f
cc_27 N_VSS_c_27_p N_VDD_c_100_n 0.00142235f
cc_28 VSS N_VDD_c_100_n 0.00104966f
cc_29 N_VSS_c_23_p N_VDD_c_104_n 3.91951e-19
cc_30 N_VSS_c_30_p N_VDD_c_104_n 8.51944e-19
cc_31 N_VSS_c_31_p N_VDD_c_104_n 3.99794e-19
cc_32 N_VSS_c_32_p N_VDD_c_107_n 3.80388e-19
cc_33 N_VSS_c_4_p N_VDD_c_107_n 3.60588e-19
cc_34 N_VSS_c_30_p N_VDD_c_107_n 0.00141604f
cc_35 N_VSS_c_31_p N_VDD_c_107_n 0.00112293f
cc_36 N_VSS_c_27_p N_VDD_c_107_n 0.00608608f
cc_37 N_VSS_c_30_p N_VDD_c_112_n 9.12964e-19
cc_38 N_VSS_c_31_p N_VDD_c_112_n 3.66936e-19
cc_39 N_VSS_c_7_p N_VDD_c_114_n 0.00116512f
cc_40 N_VSS_c_20_p N_VDD_c_115_n 9.75006e-19
cc_41 N_VSS_c_27_p N_VDD_c_116_n 9.68945e-19
cc_42 N_VSS_c_9_p N_VDD_c_117_n 3.44698e-19
cc_43 N_VSS_c_10_p N_VDD_c_117_n 7.93802e-19
cc_44 N_VSS_c_30_p N_VDD_c_119_n 3.48267e-19
cc_45 N_VSS_c_31_p N_VDD_c_119_n 8.07896e-19
cc_46 N_VSS_c_10_p N_B_c_160_n 0.00234321f
cc_47 N_VSS_c_9_p N_B_c_161_n 8.39582e-19
cc_48 N_VSS_c_10_p N_B_c_161_n 5.42695e-19
cc_49 N_VSS_c_7_p N_B_c_161_n 7.94601e-19
cc_50 N_VSS_c_10_p N_B_c_164_n 2.00604e-19
cc_51 N_VSS_c_51_p N_B_c_165_n 8.37306e-19
cc_52 N_VSS_c_9_p N_B_c_165_n 4.56568e-19
cc_53 N_VSS_c_10_p N_B_c_165_n 0.00173573f
cc_54 N_VSS_XI2.X0_S N_NET21_XI2.X0_D 3.43419e-19
cc_55 N_VSS_c_6_p N_NET21_XI2.X0_D 3.48267e-19
cc_56 N_VSS_XI1.X0_S N_NET21_XI0.X0_D 3.43419e-19
cc_57 N_VSS_c_23_p N_NET21_XI0.X0_D 3.48267e-19
cc_58 N_VSS_c_31_p N_NET21_XI4.X0_CG 7.99056e-19
cc_59 N_VSS_XI4.X0_PGD N_NET21_c_190_n 4.20799e-19
cc_60 N_VSS_XI1.X0_S N_NET21_c_191_n 3.48267e-19
cc_61 N_VSS_c_6_p N_NET21_c_191_n 8.89782e-19
cc_62 N_VSS_c_23_p N_NET21_c_191_n 5.69026e-19
cc_63 N_VSS_c_7_p N_NET21_c_191_n 2.81358e-19
cc_64 N_VSS_c_7_p N_NET21_c_195_n 2.56803e-19
cc_65 N_VSS_c_27_p N_NET21_c_195_n 2.99166e-19
cc_66 N_VSS_c_23_p N_NET21_c_197_n 9.55513e-19
cc_67 N_VSS_c_7_p N_NET21_c_197_n 2.03357e-19
cc_68 N_VSS_c_20_p N_NET21_c_197_n 9.1856e-19
cc_69 N_VSS_XI0.X0_PGD N_A_c_224_n 9.39677e-19
cc_70 N_VSS_c_3_p N_A_c_224_n 2.16729e-19
cc_71 N_VSS_XI1.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_72 N_VSS_c_23_p N_Z_XI3.X0_D 3.48267e-19
cc_73 N_VSS_XI1.X0_S N_Z_c_248_n 3.48267e-19
cc_74 N_VSS_c_23_p N_Z_c_248_n 7.85754e-19
cc_75 N_VSS_c_27_p N_Z_c_248_n 2.64173e-19
cc_76 N_VDD_c_121_p N_B_XI2.X0_CG 0.00237871f
cc_77 N_VDD_c_121_p N_B_c_169_n 0.00105622f
cc_78 N_VDD_c_80_n N_B_c_161_n 0.0025613f
cc_79 N_VDD_c_124_p N_B_c_161_n 7.31965e-19
cc_80 N_VDD_c_121_p N_B_c_161_n 5.48584e-19
cc_81 N_VDD_c_80_n N_B_c_164_n 4.9897e-19
cc_82 N_VDD_c_124_p N_B_c_164_n 4.85469e-19
cc_83 N_VDD_c_121_p N_B_c_164_n 0.00150793f
cc_84 N_VDD_c_80_n N_B_c_165_n 3.66936e-19
cc_85 N_VDD_c_121_p N_B_c_165_n 2.00604e-19
cc_86 N_VDD_XI0.X0_S N_NET21_XI0.X0_D 3.43419e-19
cc_87 N_VDD_c_90_n N_NET21_XI0.X0_D 3.72199e-19
cc_88 N_VDD_c_91_n N_NET21_XI0.X0_D 3.7884e-19
cc_89 N_VDD_c_119_n N_NET21_c_203_n 0.00250475f
cc_90 N_VDD_XI3.X0_PGD N_NET21_c_190_n 4.25379e-19
cc_91 N_VDD_XI0.X0_S N_NET21_c_191_n 3.48267e-19
cc_92 N_VDD_c_80_n N_NET21_c_191_n 4.38672e-19
cc_93 N_VDD_c_90_n N_NET21_c_191_n 7.89245e-19
cc_94 N_VDD_c_91_n N_NET21_c_191_n 5.36364e-19
cc_95 N_VDD_c_140_p N_NET21_c_195_n 3.64358e-19
cc_96 N_VDD_c_104_n N_NET21_c_195_n 6.84156e-19
cc_97 N_VDD_c_119_n N_NET21_c_195_n 4.99367e-19
cc_98 N_VDD_c_104_n N_NET21_c_212_n 4.85469e-19
cc_99 N_VDD_c_119_n N_NET21_c_212_n 0.0014909f
cc_100 N_VDD_XI2.X0_PGD N_A_c_224_n 5.10213e-19
cc_101 N_VDD_XI1.X0_PGD N_A_c_224_n 2.48727e-19
cc_102 N_VDD_XI2.X0_PGS N_A_c_228_n 6.4837e-19
cc_103 N_VDD_c_80_n N_A_c_228_n 3.16598e-19
cc_104 N_VDD_c_149_p N_A_c_230_n 8.9931e-19
cc_105 N_VDD_c_97_n N_A_c_230_n 4.91217e-19
cc_106 N_VDD_c_117_n N_A_c_230_n 0.00142365f
cc_107 N_VDD_c_97_n A 6.02732e-19
cc_108 N_VDD_c_117_n A 4.56568e-19
cc_109 N_VDD_XI4.X0_S N_Z_XI3.X0_D 3.43419e-19
cc_110 N_VDD_c_107_n N_Z_XI3.X0_D 3.7884e-19
cc_111 N_VDD_c_156_p N_Z_XI3.X0_D 3.72199e-19
cc_112 N_VDD_XI4.X0_S N_Z_c_248_n 3.48267e-19
cc_113 N_VDD_c_107_n N_Z_c_248_n 5.12447e-19
cc_114 N_VDD_c_156_p N_Z_c_248_n 7.4527e-19
cc_115 N_B_c_161_n N_NET21_c_191_n 0.00757794f
cc_116 N_B_c_164_n N_NET21_c_191_n 9.56873e-19
cc_117 N_B_c_165_n N_NET21_c_191_n 8.92526e-19
cc_118 N_B_c_160_n N_A_XI0.X0_PGS 4.5346e-19
cc_119 N_B_c_165_n N_A_XI0.X0_PGS 7.86826e-19
cc_120 N_B_c_164_n N_A_c_224_n 9.25308e-19
cc_121 N_B_c_165_n N_A_c_230_n 7.50183e-19
cc_122 N_NET21_c_191_n N_A_c_224_n 8.63036e-19
cc_123 N_NET21_c_191_n N_A_c_230_n 9.38449e-19
cc_124 N_NET21_c_195_n N_A_c_230_n 3.48267e-19
cc_125 N_NET21_c_212_n N_A_c_230_n 0.00196751f
cc_126 N_NET21_c_191_n A 0.00142917f
cc_127 N_NET21_c_195_n A 4.28721e-19
cc_128 N_NET21_c_197_n A 3.26205e-19
*
.ends
*
*
.subckt OR2_HPNW4 A B Y VDD VSS
xgate (VSS VDD B A Y) G3_OR2_N1
.ends
*
* File: G4_XNOR2_N1.pex.netlist
* Created: Wed Mar 16 10:29:55 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XNOR2_N1_VDD 2 5 9 12 16 32 35 42 43 66 68 69 70 73 75 76 79 81 85
+ 89 91 93 98 99 100 103 109 114 Vss
c113 114 Vss 0.00462632f
c114 109 Vss 0.00491723f
c115 101 Vss 8.54719e-19
c116 100 Vss 2.39889e-19
c117 99 Vss 3.56526e-19
c118 98 Vss 0.0049606f
c119 93 Vss 0.00247173f
c120 91 Vss 0.0107823f
c121 89 Vss 0.00155915f
c122 85 Vss 3.94646e-19
c123 81 Vss 0.00431979f
c124 79 Vss 0.00104496f
c125 76 Vss 8.67334e-19
c126 75 Vss 0.00219831f
c127 73 Vss 0.00159894f
c128 70 Vss 8.63261e-19
c129 69 Vss 0.00531705f
c130 68 Vss 0.00645016f
c131 66 Vss 0.00203422f
c132 43 Vss 0.0336444f
c133 42 Vss 0.0994765f
c134 35 Vss 7.78608e-20
c135 33 Vss 0.0348624f
c136 32 Vss 0.0999592f
c137 16 Vss 0.00272748f
c138 12 Vss 0.00264503f
c139 9 Vss 0.165252f
c140 5 Vss 0.165777f
c141 2 Vss 0.00272748f
r142 98 103 0.326018
r143 97 98 4.16786
r144 93 97 0.655813
r145 93 95 1.82344
r146 92 101 0.494161
r147 91 103 0.326018
r148 91 92 13.0037
r149 87 101 0.128424
r150 87 89 4.83471
r151 85 114 1.16709
r152 83 85 2.16729
r153 82 100 0.494161
r154 81 101 0.494161
r155 81 82 7.46046
r156 79 109 1.16709
r157 77 100 0.128424
r158 77 79 2.16729
r159 75 100 0.494161
r160 75 76 4.37625
r161 71 99 0.0828784
r162 71 73 1.82344
r163 69 83 0.652036
r164 69 70 10.1279
r165 68 76 0.652036
r166 67 99 0.551426
r167 67 68 12.1701
r168 66 99 0.551426
r169 65 70 0.652036
r170 65 66 4.16786
r171 45 114 0.238214
r172 43 45 1.45875
r173 42 46 0.652036
r174 42 45 1.45875
r175 39 43 0.652036
r176 35 109 0.238214
r177 33 35 1.45875
r178 32 36 0.652036
r179 32 35 1.45875
r180 29 33 0.652036
r181 16 95 1.16709
r182 12 89 1.16709
r183 9 46 2.5674
r184 9 39 2.5674
r185 5 36 2.5674
r186 5 29 2.5674
r187 2 73 1.16709
.ends

.subckt PM_G4_XNOR2_N1_VSS 3 6 8 11 16 32 33 42 43 66 71 76 81 87 96 101 114 116
+ 117 118 123 124 129 137 142 143 144 146 Vss
c99 144 Vss 3.75522e-19
c100 143 Vss 3.21033e-19
c101 142 Vss 0.00224529f
c102 141 Vss 0.0013489f
c103 137 Vss 0.00215359f
c104 129 Vss 0.0112621f
c105 124 Vss 8.17415e-19
c106 123 Vss 0.00403195f
c107 118 Vss 8.39382e-19
c108 117 Vss 0.00163605f
c109 116 Vss 0.00144702f
c110 114 Vss 0.00415033f
c111 101 Vss 0.00449981f
c112 96 Vss 0.00516182f
c113 87 Vss 7.10513e-22
c114 81 Vss 0.00255515f
c115 76 Vss 9.53239e-19
c116 71 Vss 0.00133653f
c117 66 Vss 0.00143917f
c118 43 Vss 0.033325f
c119 42 Vss 0.0990666f
c120 33 Vss 0.0336725f
c121 32 Vss 0.0976281f
c122 16 Vss 0.00213567f
c123 11 Vss 0.165384f
c124 8 Vss 0.00163738f
c125 6 Vss 0.00213969f
c126 3 Vss 0.166856f
r127 141 146 0.326018
r128 141 142 4.16786
r129 137 142 0.655813
r130 130 144 0.494161
r131 129 146 0.326018
r132 125 144 0.128424
r133 123 133 0.652036
r134 123 124 10.1279
r135 119 143 0.0828784
r136 117 144 0.494161
r137 117 118 4.37625
r138 116 124 0.652036
r139 115 143 0.551426
r140 115 116 4.16786
r141 114 143 0.551426
r142 113 118 0.652036
r143 113 114 12.1701
r144 87 137 1.82344
r145 81 129 13.5872
r146 81 130 8.04396
r147 81 84 5.37654
r148 76 101 1.16709
r149 76 133 2.16729
r150 71 96 1.16709
r151 71 125 2.16729
r152 66 119 1.82344
r153 45 101 0.238214
r154 43 45 1.45875
r155 42 46 0.652036
r156 42 45 1.45875
r157 39 43 0.652036
r158 35 96 0.238214
r159 33 35 1.45875
r160 32 36 0.652036
r161 32 35 1.45875
r162 29 33 0.652036
r163 16 87 1.16709
r164 11 46 2.5674
r165 11 39 2.5674
r166 8 84 1.16709
r167 6 66 1.16709
r168 3 36 2.5674
r169 3 29 2.5674
.ends

.subckt PM_G4_XNOR2_N1_A 2 4 7 10 18 21 24 28 39 48 51 54 57 62 67 72 77 85 Vss
c60 85 Vss 9.00557e-19
c61 77 Vss 0.00241581f
c62 72 Vss 0.00594049f
c63 67 Vss 0.00360869f
c64 62 Vss 0.00199403f
c65 57 Vss 0.00406361f
c66 51 Vss 8.38354e-19
c67 48 Vss 0.124108f
c68 43 Vss 0.0295947f
c69 39 Vss 4.97883e-20
c70 28 Vss 0.152592f
c71 24 Vss 2.44824e-19
c72 21 Vss 0.169386f
c73 18 Vss 0.0714048f
c74 16 Vss 0.0247918f
c75 10 Vss 0.0674191f
c76 7 Vss 0.219196f
c77 4 Vss 0.08397f
r78 81 85 0.653045
r79 62 77 1.16709
r80 62 85 4.9014
r81 57 72 1.16709
r82 57 81 7.87725
r83 51 67 1.16709
r84 51 54 0.0416786
r85 47 72 0.262036
r86 47 48 2.334
r87 44 47 2.20433
r88 39 77 0.404964
r89 33 48 0.00605528
r90 31 44 0.00605528
r91 29 43 0.494161
r92 28 30 0.652036
r93 28 29 4.84305
r94 25 43 0.128424
r95 24 67 0.0476429
r96 22 24 0.326018
r97 22 24 0.1167
r98 21 43 0.494161
r99 21 24 6.7686
r100 18 67 0.357321
r101 16 24 0.326018
r102 16 18 0.40845
r103 10 39 2.04225
r104 7 33 2.5674
r105 7 31 2.5674
r106 7 30 2.5674
r107 4 25 2.5674
r108 2 18 2.15895
.ends

.subckt PM_G4_XNOR2_N1_NET1 2 7 10 31 35 44 49 58 66 Vss
c38 66 Vss 6.40075e-20
c39 58 Vss 0.00598766f
c40 49 Vss 0.00482775f
c41 44 Vss 0.00129308f
c42 35 Vss 0.126399f
c43 31 Vss 0.128923f
c44 10 Vss 0.135805f
c45 7 Vss 0.297098f
c46 2 Vss 0.0015894f
r47 62 66 0.653045
r48 49 58 1.16709
r49 49 66 12.9148
r50 44 62 2.08393
r51 33 35 1.45875
r52 30 58 0.262036
r53 30 31 2.20433
r54 27 30 2.334
r55 25 35 0.259088
r56 24 31 0.00605528
r57 21 33 0.259088
r58 18 27 0.00605528
r59 10 21 4.25955
r60 7 25 5.30985
r61 7 24 2.5674
r62 7 18 2.5674
r63 2 44 1.16709
.ends

.subckt PM_G4_XNOR2_N1_NET2 2 6 9 21 22 33 42 47 56 74 Vss
c50 74 Vss 3.88292e-19
c51 56 Vss 0.00473316f
c52 47 Vss 0.00694068f
c53 42 Vss 0.00195908f
c54 33 Vss 0.123617f
c55 22 Vss 0.0344905f
c56 21 Vss 0.177827f
c57 9 Vss 0.362751f
c58 6 Vss 0.0802803f
c59 2 Vss 0.0015894f
r60 70 74 0.660011
r61 47 56 1.16709
r62 47 74 11.3611
r63 42 70 1.95889
r64 32 56 0.262036
r65 32 33 2.26917
r66 29 32 2.26917
r67 26 33 0.00605528
r68 24 29 0.00605528
r69 21 23 0.652036
r70 21 22 4.84305
r71 18 22 0.652036
r72 9 26 2.5674
r73 9 24 2.5674
r74 9 23 7.4688
r75 6 18 2.5674
r76 2 42 1.16709
.ends

.subckt PM_G4_XNOR2_N1_B 2 4 7 10 19 20 28 33 37 38 48 52 55 58 61 Vss
c37 61 Vss 0.0280185f
c38 55 Vss 9.41292e-19
c39 52 Vss 0.134888f
c40 48 Vss 0.0597924f
c41 38 Vss 0.0333789f
c42 37 Vss 0.090068f
c43 33 Vss 0.0345164f
c44 28 Vss 0.0897381f
c45 20 Vss 0.0343755f
c46 19 Vss 0.169386f
c47 10 Vss 0.155214f
c48 7 Vss 0.216f
c49 4 Vss 0.0714224f
c50 2 Vss 0.0847975f
r51 55 61 1.16709
r52 55 58 0.166714
r53 50 52 4.53833
r54 47 48 1.167
r55 42 52 0.00605528
r56 37 39 0.652036
r57 37 38 2.04225
r58 35 48 0.0685365
r59 34 50 0.00605528
r60 33 38 0.652036
r61 32 47 0.0685365
r62 32 33 1.2837
r63 31 61 0.181909
r64 29 61 0.494161
r65 29 31 0.1167
r66 28 47 0.5835
r67 28 31 3.55935
r68 23 61 0.128424
r69 23 61 0.40845
r70 22 61 0.181909
r71 20 22 6.7686
r72 19 61 0.494161
r73 19 22 0.1167
r74 16 20 0.652036
r75 10 39 5.0181
r76 7 42 2.5674
r77 7 35 2.5674
r78 7 34 2.5674
r79 4 61 2.15895
r80 2 16 2.5674
.ends

.subckt PM_G4_XNOR2_N1_Z 2 4 30 33 Vss
c27 30 Vss 0.00253242f
c28 4 Vss 0.00249005f
c29 2 Vss 0.00153036f
r30 33 35 2.9175
r31 30 33 5.08479
r32 4 35 1.16709
r33 2 30 1.16709
.ends

.subckt G4_XNOR2_N1  VDD VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI1.X0 N_NET1_XI1.X0_D N_VSS_XI1.X0_PGD N_B_XI1.X0_CG N_VSS_XI1.X0_PGD
+ N_VDD_XI1.X0_S TIGFET_HPNW4
XI9.X0 N_NET2_XI9.X0_D N_VDD_XI9.X0_PGD N_A_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI10.X0 N_NET1_XI1.X0_D N_VDD_XI10.X0_PGD N_B_XI10.X0_CG N_VDD_XI10.X0_PGD
+ N_VSS_XI10.X0_S TIGFET_HPNW4
XI3.X0 N_NET2_XI9.X0_D N_VSS_XI3.X0_PGD N_A_XI3.X0_CG N_VSS_XI3.X0_PGD
+ N_VDD_XI3.X0_S TIGFET_HPNW4
XI5.X0 N_Z_XI5.X0_D N_B_XI5.X0_PGD N_NET2_XI5.X0_CG N_B_XI5.X0_PGD
+ N_VSS_XI10.X0_S TIGFET_HPNW4
XI8.X0 N_Z_XI8.X0_D N_A_XI8.X0_PGD N_B_XI8.X0_CG N_A_XI8.X0_PGD N_VDD_XI3.X0_S
+ TIGFET_HPNW4
XI11.X0 N_Z_XI5.X0_D N_NET1_XI11.X0_PGD N_A_XI11.X0_CG N_NET1_XI11.X0_PGD
+ N_VSS_XI11.X0_S TIGFET_HPNW4
XI7.X0 N_Z_XI8.X0_D N_NET2_XI7.X0_PGD N_NET1_XI7.X0_CG N_NET2_XI7.X0_PGD
+ N_VDD_XI7.X0_S TIGFET_HPNW4
*
x_PM_G4_XNOR2_N1_VDD N_VDD_XI1.X0_S N_VDD_XI9.X0_PGD N_VDD_XI10.X0_PGD
+ N_VDD_XI3.X0_S N_VDD_XI7.X0_S N_VDD_c_11_p N_VDD_c_58_p N_VDD_c_26_p
+ N_VDD_c_8_p N_VDD_c_17_p N_VDD_c_14_p N_VDD_c_9_p N_VDD_c_45_p N_VDD_c_3_p
+ N_VDD_c_16_p N_VDD_c_49_p N_VDD_c_21_p N_VDD_c_12_p N_VDD_c_19_p N_VDD_c_4_p
+ N_VDD_c_60_p N_VDD_c_7_p N_VDD_c_90_p N_VDD_c_42_p N_VDD_c_48_p VDD
+ N_VDD_c_24_p N_VDD_c_20_p Vss PM_G4_XNOR2_N1_VDD
x_PM_G4_XNOR2_N1_VSS N_VSS_XI1.X0_PGD N_VSS_XI9.X0_S N_VSS_XI10.X0_S
+ N_VSS_XI3.X0_PGD N_VSS_XI11.X0_S N_VSS_c_121_n N_VSS_c_123_n N_VSS_c_172_p
+ N_VSS_c_124_n N_VSS_c_126_n N_VSS_c_130_n N_VSS_c_134_n N_VSS_c_138_n
+ N_VSS_c_143_n N_VSS_c_145_n N_VSS_c_149_n N_VSS_c_153_n N_VSS_c_156_n
+ N_VSS_c_157_n N_VSS_c_158_n N_VSS_c_159_n N_VSS_c_162_n N_VSS_c_163_n
+ N_VSS_c_164_n N_VSS_c_185_p N_VSS_c_165_n N_VSS_c_166_n VSS Vss
+ PM_G4_XNOR2_N1_VSS
x_PM_G4_XNOR2_N1_A N_A_XI9.X0_CG N_A_XI3.X0_CG N_A_XI8.X0_PGD N_A_XI11.X0_CG
+ N_A_c_214_n N_A_c_215_n N_A_c_217_n N_A_c_218_n N_A_c_249_p N_A_c_219_n
+ N_A_c_220_n A N_A_c_223_n N_A_c_225_n N_A_c_226_n N_A_c_229_n N_A_c_244_p
+ N_A_c_242_n Vss PM_G4_XNOR2_N1_A
x_PM_G4_XNOR2_N1_NET1 N_NET1_XI1.X0_D N_NET1_XI11.X0_PGD N_NET1_XI7.X0_CG
+ N_NET1_c_309_p N_NET1_c_293_n N_NET1_c_276_n N_NET1_c_279_n N_NET1_c_296_n
+ N_NET1_c_280_n Vss PM_G4_XNOR2_N1_NET1
x_PM_G4_XNOR2_N1_NET2 N_NET2_XI9.X0_D N_NET2_XI5.X0_CG N_NET2_XI7.X0_PGD
+ N_NET2_c_336_n N_NET2_c_356_p N_NET2_c_314_n N_NET2_c_315_n N_NET2_c_318_n
+ N_NET2_c_322_n N_NET2_c_324_n Vss PM_G4_XNOR2_N1_NET2
x_PM_G4_XNOR2_N1_B N_B_XI1.X0_CG N_B_XI10.X0_CG N_B_XI5.X0_PGD N_B_XI8.X0_CG
+ N_B_c_363_n N_B_c_382_n N_B_c_365_n N_B_c_392_n N_B_c_388_n N_B_c_384_n
+ N_B_c_395_n N_B_c_366_n N_B_c_367_n B N_B_c_369_n Vss PM_G4_XNOR2_N1_B
x_PM_G4_XNOR2_N1_Z N_Z_XI5.X0_D N_Z_XI8.X0_D N_Z_c_403_n Z Vss PM_G4_XNOR2_N1_Z
cc_1 N_VDD_XI9.X0_PGD N_VSS_XI1.X0_PGD 2.96813e-19
cc_2 N_VDD_XI10.X0_PGD N_VSS_XI1.X0_PGD 0.00168295f
cc_3 N_VDD_c_3_p N_VSS_XI9.X0_S 2.15082e-19
cc_4 N_VDD_c_4_p N_VSS_XI10.X0_S 2.35318e-19
cc_5 N_VDD_XI9.X0_PGD N_VSS_XI3.X0_PGD 0.00167677f
cc_6 N_VDD_c_4_p N_VSS_XI3.X0_PGD 2.68479e-19
cc_7 N_VDD_c_7_p N_VSS_XI11.X0_S 2.15082e-19
cc_8 N_VDD_c_8_p N_VSS_c_121_n 0.00168295f
cc_9 N_VDD_c_9_p N_VSS_c_121_n 3.60588e-19
cc_10 N_VDD_c_9_p N_VSS_c_123_n 3.60588e-19
cc_11 N_VDD_c_11_p N_VSS_c_124_n 0.00167677f
cc_12 N_VDD_c_12_p N_VSS_c_124_n 3.60588e-19
cc_13 N_VDD_XI1.X0_S N_VSS_c_126_n 2.15082e-19
cc_14 N_VDD_c_14_p N_VSS_c_126_n 0.00187494f
cc_15 N_VDD_c_3_p N_VSS_c_126_n 8.9077e-19
cc_16 N_VDD_c_16_p N_VSS_c_126_n 5.16845e-19
cc_17 N_VDD_c_17_p N_VSS_c_130_n 4.43871e-19
cc_18 N_VDD_c_9_p N_VSS_c_130_n 0.00141228f
cc_19 N_VDD_c_19_p N_VSS_c_130_n 8.52111e-19
cc_20 N_VDD_c_20_p N_VSS_c_130_n 3.48267e-19
cc_21 N_VDD_c_21_p N_VSS_c_134_n 9.21268e-19
cc_22 N_VDD_c_12_p N_VSS_c_134_n 0.00141228f
cc_23 N_VDD_c_4_p N_VSS_c_134_n 0.00225084f
cc_24 N_VDD_c_24_p N_VSS_c_134_n 3.48267e-19
cc_25 N_VDD_XI3.X0_S N_VSS_c_138_n 2.35318e-19
cc_26 N_VDD_c_26_p N_VSS_c_138_n 2.72094e-19
cc_27 N_VDD_c_9_p N_VSS_c_138_n 0.00534617f
cc_28 N_VDD_c_4_p N_VSS_c_138_n 4.25159e-19
cc_29 N_VDD_c_20_p N_VSS_c_138_n 9.58524e-19
cc_30 N_VDD_XI7.X0_S N_VSS_c_143_n 2.15082e-19
cc_31 N_VDD_c_7_p N_VSS_c_143_n 3.16299e-19
cc_32 N_VDD_c_17_p N_VSS_c_145_n 3.66936e-19
cc_33 N_VDD_c_9_p N_VSS_c_145_n 0.00112249f
cc_34 N_VDD_c_19_p N_VSS_c_145_n 3.99794e-19
cc_35 N_VDD_c_20_p N_VSS_c_145_n 8.03027e-19
cc_36 N_VDD_c_21_p N_VSS_c_149_n 3.82294e-19
cc_37 N_VDD_c_12_p N_VSS_c_149_n 0.00112249f
cc_38 N_VDD_c_4_p N_VSS_c_149_n 9.55322e-19
cc_39 N_VDD_c_24_p N_VSS_c_149_n 8.0279e-19
cc_40 N_VDD_c_17_p N_VSS_c_153_n 0.00287902f
cc_41 N_VDD_c_14_p N_VSS_c_153_n 0.0057117f
cc_42 N_VDD_c_42_p N_VSS_c_153_n 0.0010706f
cc_43 N_VDD_c_14_p N_VSS_c_156_n 0.00304013f
cc_44 N_VDD_c_9_p N_VSS_c_157_n 0.00342836f
cc_45 N_VDD_c_45_p N_VSS_c_158_n 0.00107429f
cc_46 N_VDD_c_16_p N_VSS_c_159_n 0.00352516f
cc_47 N_VDD_c_12_p N_VSS_c_159_n 0.0060405f
cc_48 N_VDD_c_48_p N_VSS_c_159_n 0.00101104f
cc_49 N_VDD_c_49_p N_VSS_c_162_n 0.00105833f
cc_50 N_VDD_c_9_p N_VSS_c_163_n 0.00458401f
cc_51 N_VDD_c_7_p N_VSS_c_164_n 0.00135143f
cc_52 N_VDD_c_14_p N_VSS_c_165_n 7.88896e-19
cc_53 N_VDD_c_9_p N_VSS_c_166_n 7.74609e-19
cc_54 N_VDD_c_4_p N_A_XI8.X0_PGD 2.51969e-19
cc_55 N_VDD_c_24_p N_A_c_214_n 0.00237738f
cc_56 N_VDD_XI9.X0_PGD N_A_c_215_n 4.04053e-19
cc_57 N_VDD_XI10.X0_PGD N_A_c_215_n 2.40582e-19
cc_58 N_VDD_c_58_p N_A_c_217_n 9.54306e-19
cc_59 N_VDD_XI10.X0_PGD N_A_c_218_n 2.40582e-19
cc_60 N_VDD_c_60_p N_A_c_219_n 5.838e-19
cc_61 N_VDD_c_14_p N_A_c_220_n 5.24876e-19
cc_62 N_VDD_c_21_p N_A_c_220_n 6.41525e-19
cc_63 N_VDD_c_24_p N_A_c_220_n 4.56568e-19
cc_64 N_VDD_c_4_p N_A_c_223_n 0.00237851f
cc_65 N_VDD_c_60_p N_A_c_223_n 0.00200281f
cc_66 N_VDD_c_60_p N_A_c_225_n 8.17097e-19
cc_67 N_VDD_c_14_p N_A_c_226_n 6.27972e-19
cc_68 N_VDD_c_21_p N_A_c_226_n 4.85469e-19
cc_69 N_VDD_c_24_p N_A_c_226_n 6.1245e-19
cc_70 N_VDD_c_4_p N_A_c_229_n 9.84209e-19
cc_71 N_VDD_c_60_p N_A_c_229_n 2.37583e-19
cc_72 N_VDD_XI1.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_73 N_VDD_c_9_p N_NET1_XI1.X0_D 3.7884e-19
cc_74 N_VDD_c_3_p N_NET1_XI1.X0_D 3.72199e-19
cc_75 N_VDD_XI1.X0_S N_NET1_c_276_n 3.48267e-19
cc_76 N_VDD_c_9_p N_NET1_c_276_n 4.58491e-19
cc_77 N_VDD_c_3_p N_NET1_c_276_n 5.226e-19
cc_78 N_VDD_c_19_p N_NET1_c_279_n 0.00121121f
cc_79 N_VDD_c_9_p N_NET1_c_280_n 3.78572e-19
cc_80 N_VDD_XI3.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_81 N_VDD_c_12_p N_NET2_XI9.X0_D 3.7884e-19
cc_82 N_VDD_c_4_p N_NET2_XI9.X0_D 3.48267e-19
cc_83 N_VDD_c_60_p N_NET2_c_314_n 8.01015e-19
cc_84 N_VDD_XI3.X0_S N_NET2_c_315_n 3.48267e-19
cc_85 N_VDD_c_12_p N_NET2_c_315_n 4.58491e-19
cc_86 N_VDD_c_4_p N_NET2_c_315_n 8.45449e-19
cc_87 N_VDD_c_12_p N_NET2_c_318_n 3.29894e-19
cc_88 N_VDD_c_4_p N_NET2_c_318_n 8.51778e-19
cc_89 N_VDD_c_60_p N_NET2_c_318_n 0.00334727f
cc_90 N_VDD_c_90_p N_NET2_c_318_n 7.7731e-19
cc_91 N_VDD_c_60_p N_NET2_c_322_n 2.33029e-19
cc_92 N_VDD_c_90_p N_NET2_c_322_n 3.66936e-19
cc_93 N_VDD_c_21_p N_NET2_c_324_n 3.10284e-19
cc_94 N_VDD_c_20_p N_B_XI10.X0_CG 0.00237871f
cc_95 N_VDD_XI10.X0_PGD N_B_XI5.X0_PGD 0.00176522f
cc_96 N_VDD_XI9.X0_PGD N_B_c_363_n 2.40582e-19
cc_97 N_VDD_XI10.X0_PGD N_B_c_363_n 4.04053e-19
cc_98 N_VDD_XI10.X0_PGD N_B_c_365_n 4.05198e-19
cc_99 N_VDD_c_26_p N_B_c_366_n 0.00154836f
cc_100 N_VDD_c_19_p N_B_c_367_n 5.50671e-19
cc_101 N_VDD_c_20_p N_B_c_367_n 8.9014e-19
cc_102 N_VDD_c_19_p N_B_c_369_n 4.73723e-19
cc_103 N_VDD_c_20_p N_B_c_369_n 0.0014909f
cc_104 N_VDD_XI3.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_105 N_VDD_XI7.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_106 N_VDD_c_4_p N_Z_XI8.X0_D 3.48267e-19
cc_107 N_VDD_c_60_p N_Z_XI8.X0_D 3.7884e-19
cc_108 N_VDD_c_7_p N_Z_XI8.X0_D 3.72199e-19
cc_109 N_VDD_XI3.X0_S N_Z_c_403_n 3.48267e-19
cc_110 N_VDD_XI7.X0_S N_Z_c_403_n 3.48267e-19
cc_111 N_VDD_c_4_p N_Z_c_403_n 5.21254e-19
cc_112 N_VDD_c_60_p N_Z_c_403_n 6.55718e-19
cc_113 N_VDD_c_7_p N_Z_c_403_n 8.25922e-19
cc_114 N_VSS_c_149_n N_A_XI3.X0_CG 9.02944e-19
cc_115 N_VSS_XI3.X0_PGD N_A_XI8.X0_PGD 0.00150976f
cc_116 N_VSS_XI1.X0_PGD N_A_c_215_n 2.40582e-19
cc_117 N_VSS_XI3.X0_PGD N_A_c_215_n 3.99472e-19
cc_118 N_VSS_XI3.X0_PGD N_A_c_218_n 4.05198e-19
cc_119 N_VSS_c_172_p N_A_c_219_n 0.00150976f
cc_120 N_VSS_c_134_n N_A_c_223_n 4.12959e-19
cc_121 N_VSS_c_153_n N_A_c_223_n 3.96361e-19
cc_122 N_VSS_c_163_n N_A_c_225_n 2.41875e-19
cc_123 N_VSS_c_145_n N_A_c_226_n 4.65658e-19
cc_124 N_VSS_c_149_n N_A_c_229_n 8.90609e-19
cc_125 N_VSS_c_163_n N_A_c_242_n 3.10545e-19
cc_126 N_VSS_XI10.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_127 N_VSS_c_138_n N_NET1_XI1.X0_D 3.48267e-19
cc_128 N_VSS_XI10.X0_S N_NET1_c_276_n 3.48267e-19
cc_129 N_VSS_c_138_n N_NET1_c_276_n 0.0012813f
cc_130 N_VSS_c_138_n N_NET1_c_279_n 0.00174104f
cc_131 N_VSS_c_163_n N_NET1_c_279_n 5.89244e-19
cc_132 N_VSS_c_185_p N_NET1_c_279_n 0.00121599f
cc_133 N_VSS_c_130_n N_NET1_c_280_n 0.00206231f
cc_134 N_VSS_c_153_n N_NET1_c_280_n 9.32604e-19
cc_135 N_VSS_c_163_n N_NET1_c_280_n 0.0214545f
cc_136 N_VSS_XI9.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_137 N_VSS_c_126_n N_NET2_XI9.X0_D 3.48267e-19
cc_138 N_VSS_XI9.X0_S N_NET2_c_315_n 3.48267e-19
cc_139 N_VSS_c_126_n N_NET2_c_315_n 0.00108327f
cc_140 N_VSS_c_159_n N_NET2_c_315_n 3.31434e-19
cc_141 N_VSS_c_134_n N_NET2_c_318_n 0.00143089f
cc_142 N_VSS_c_156_n N_NET2_c_324_n 3.36104e-19
cc_143 N_VSS_c_159_n N_NET2_c_324_n 6.48614e-19
cc_144 N_VSS_c_145_n N_B_XI1.X0_CG 9.02944e-19
cc_145 N_VSS_XI1.X0_PGD N_B_c_363_n 3.99472e-19
cc_146 N_VSS_XI3.X0_PGD N_B_c_363_n 2.40582e-19
cc_147 N_VSS_XI3.X0_PGD N_B_c_365_n 2.40582e-19
cc_148 N_VSS_c_138_n N_B_c_366_n 2.8419e-19
cc_149 N_VSS_c_149_n N_B_c_367_n 2.07877e-19
cc_150 N_VSS_c_153_n N_B_c_367_n 2.27769e-19
cc_151 N_VSS_c_149_n N_B_c_369_n 7.33679e-19
cc_152 N_VSS_XI10.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_153 N_VSS_XI11.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_154 N_VSS_c_138_n N_Z_XI5.X0_D 3.48267e-19
cc_155 N_VSS_c_143_n N_Z_XI5.X0_D 3.48267e-19
cc_156 N_VSS_XI10.X0_S N_Z_c_403_n 3.48267e-19
cc_157 N_VSS_XI11.X0_S N_Z_c_403_n 3.48267e-19
cc_158 N_VSS_c_138_n N_Z_c_403_n 8.61925e-19
cc_159 N_VSS_c_143_n N_Z_c_403_n 5.69026e-19
cc_160 N_A_XI11.X0_CG N_NET1_XI11.X0_PGD 4.5346e-19
cc_161 N_A_c_244_p N_NET1_XI11.X0_PGD 0.00151381f
cc_162 N_A_c_244_p N_NET1_c_293_n 0.00157635f
cc_163 N_A_c_225_n N_NET1_c_279_n 0.00310276f
cc_164 N_A_c_242_n N_NET1_c_279_n 0.00205512f
cc_165 N_A_XI11.X0_CG N_NET1_c_296_n 0.00234108f
cc_166 N_A_c_249_p N_NET1_c_296_n 0.00101616f
cc_167 N_A_c_244_p N_NET1_c_296_n 0.00161406f
cc_168 N_A_XI8.X0_PGD N_NET2_XI7.X0_PGD 0.00160287f
cc_169 N_A_c_218_n N_NET2_XI7.X0_PGD 3.14428e-19
cc_170 N_A_c_244_p N_NET2_XI7.X0_PGD 5.68075e-19
cc_171 N_A_XI8.X0_PGD N_NET2_c_336_n 4.60549e-19
cc_172 N_A_c_219_n N_NET2_c_314_n 0.00160287f
cc_173 N_A_c_223_n N_NET2_c_315_n 7.37727e-19
cc_174 N_A_c_223_n N_NET2_c_318_n 0.00205074f
cc_175 N_A_c_225_n N_NET2_c_318_n 0.0018485f
cc_176 N_A_c_229_n N_NET2_c_318_n 3.44698e-19
cc_177 N_A_c_223_n N_NET2_c_322_n 3.44698e-19
cc_178 N_A_c_229_n N_NET2_c_322_n 9.07485e-19
cc_179 N_A_c_244_p N_NET2_c_322_n 3.98239e-19
cc_180 N_A_c_218_n N_B_XI8.X0_CG 0.003858f
cc_181 N_A_c_229_n N_B_XI8.X0_CG 0.00111269f
cc_182 N_A_c_215_n N_B_c_363_n 0.00575421f
cc_183 N_A_c_226_n N_B_c_382_n 4.09767e-19
cc_184 N_A_c_218_n N_B_c_365_n 0.00308843f
cc_185 N_A_c_218_n N_B_c_384_n 0.00362155f
cc_186 N_A_c_215_n N_B_c_369_n 6.77269e-19
cc_187 N_A_c_223_n N_Z_c_403_n 0.00321233f
cc_188 N_A_c_225_n N_Z_c_403_n 0.0025035f
cc_189 N_A_c_244_p N_Z_c_403_n 8.50872e-19
cc_190 N_NET1_c_276_n N_NET2_XI9.X0_D 2.15082e-19
cc_191 N_NET1_XI11.X0_PGD N_NET2_XI5.X0_CG 2.62058e-19
cc_192 N_NET1_c_293_n N_NET2_XI7.X0_PGD 0.00832016f
cc_193 N_NET1_XI11.X0_PGD N_NET2_c_336_n 0.00416722f
cc_194 N_NET1_XI1.X0_D N_NET2_c_315_n 2.15082e-19
cc_195 N_NET1_c_279_n N_NET2_c_318_n 0.00142494f
cc_196 N_NET1_XI7.X0_CG N_NET2_c_322_n 0.00102831f
cc_197 N_NET1_XI11.X0_PGD N_B_XI5.X0_PGD 0.00188492f
cc_198 N_NET1_XI7.X0_CG N_B_XI8.X0_CG 2.60667e-19
cc_199 N_NET1_c_293_n N_B_c_388_n 2.60667e-19
cc_200 N_NET1_c_309_p N_B_c_366_n 0.00165894f
cc_201 N_NET1_c_279_n N_Z_c_403_n 3.02205e-19
cc_202 N_NET2_XI5.X0_CG N_B_XI5.X0_PGD 0.0019183f
cc_203 N_NET2_c_336_n N_B_XI5.X0_PGD 0.00161994f
cc_204 N_NET2_XI7.X0_PGD N_B_c_392_n 3.1641e-19
cc_205 N_NET2_XI7.X0_PGD N_B_c_388_n 0.00313953f
cc_206 N_NET2_c_356_p N_B_c_388_n 0.00172424f
cc_207 N_NET2_c_356_p N_B_c_395_n 0.0019183f
cc_208 N_NET2_XI7.X0_PGD N_Z_c_403_n 0.00115814f
cc_209 N_NET2_c_336_n N_Z_c_403_n 5.21666e-19
cc_210 N_NET2_c_318_n N_Z_c_403_n 2.80086e-19
cc_211 N_B_c_388_n N_Z_c_403_n 8.84927e-19
cc_212 N_B_c_367_n N_Z_c_403_n 3.17615e-19
*
.ends
*
*
.subckt XNOR2_HPNW4 A B Y VDD VSS
xgate (VDD VSS A B Y) G4_XNOR2_N1
.ends
*
* File: G5_XNOR3_N1.pex.netlist
* Created: Fri Mar 25 15:42:00 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XNOR3_N1_VDD 2 5 9 12 14 17 34 35 44 45 54 55 77 79 80 81 84 86 90
+ 93 96 98 102 104 108 112 114 116 118 119 125 134 139 Vss
c122 139 Vss 0.00481852f
c123 134 Vss 0.00580927f
c124 125 Vss 0.00558883f
c125 119 Vss 2.39889e-19
c126 118 Vss 4.91159e-19
c127 117 Vss 4.14624e-19
c128 114 Vss 3.56526e-19
c129 112 Vss 0.00104518f
c130 108 Vss 3.94646e-19
c131 104 Vss 0.00602085f
c132 102 Vss 0.00109141f
c133 98 Vss 0.00553212f
c134 96 Vss 0.0016276f
c135 93 Vss 0.00243759f
c136 90 Vss 0.00352468f
c137 86 Vss 0.00659816f
c138 84 Vss 0.0015095f
c139 81 Vss 8.67152e-19
c140 80 Vss 0.00945954f
c141 79 Vss 0.00914208f
c142 77 Vss 0.00176824f
c143 57 Vss 5.45153e-20
c144 55 Vss 0.0336444f
c145 54 Vss 0.0988545f
c146 45 Vss 0.0346156f
c147 44 Vss 0.1003f
c148 35 Vss 0.0346129f
c149 34 Vss 0.0990563f
c150 17 Vss 0.165098f
c151 14 Vss 0.00210084f
c152 12 Vss 0.00231756f
c153 9 Vss 0.16518f
c154 5 Vss 0.165156f
c155 2 Vss 0.00208065f
r156 110 112 4.83471
r157 108 139 1.16709
r158 106 108 2.16729
r159 105 119 0.494161
r160 104 110 0.652036
r161 104 105 7.46046
r162 102 134 1.16709
r163 100 119 0.128424
r164 100 102 2.16729
r165 99 118 0.494161
r166 98 106 0.652036
r167 98 99 10.3363
r168 94 117 0.0828784
r169 94 96 2.00578
r170 93 118 0.128424
r171 92 117 0.551426
r172 92 93 4.16786
r173 90 125 1.16709
r174 88 117 0.551426
r175 88 90 5.835
r176 87 116 0.326018
r177 86 118 0.494161
r178 86 87 10.1279
r179 82 114 0.0828784
r180 82 84 1.82344
r181 80 119 0.494161
r182 80 81 15.8795
r183 79 116 0.326018
r184 78 114 0.551426
r185 78 79 13.3371
r186 77 114 0.551426
r187 76 81 0.652036
r188 76 77 4.16786
r189 57 139 0.238214
r190 55 57 1.45875
r191 54 58 0.652036
r192 54 57 1.45875
r193 51 55 0.652036
r194 47 134 0.238214
r195 45 47 1.45875
r196 44 48 0.652036
r197 44 47 1.45875
r198 41 45 0.652036
r199 37 125 0.238214
r200 35 37 1.45875
r201 34 38 0.652036
r202 34 37 1.45875
r203 31 35 0.652036
r204 17 58 2.5674
r205 17 51 2.5674
r206 14 112 1.16709
r207 12 96 1.16709
r208 9 48 2.5674
r209 9 41 2.5674
r210 5 38 2.5674
r211 5 31 2.5674
r212 2 84 1.16709
.ends

.subckt PM_G5_XNOR3_N1_C 2 4 6 8 17 20 23 40 43 47 52 57 62 85 87 93 98 Vss
c60 98 Vss 8.02961e-19
c61 93 Vss 6.27504e-19
c62 87 Vss 0.0049214f
c63 85 Vss 0.00877979f
c64 62 Vss 0.00258187f
c65 57 Vss 0.00458232f
c66 52 Vss 0.00201471f
c67 47 Vss 4.03464e-19
c68 43 Vss 3.73849e-19
c69 40 Vss 5.60764e-19
c70 23 Vss 1.05295e-19
c71 20 Vss 0.220565f
c72 17 Vss 0.0715834f
c73 15 Vss 0.0247918f
c74 8 Vss 0.00236553f
c75 4 Vss 0.0826049f
r76 88 98 0.0685365
r77 87 89 0.652036
r78 87 88 10.3363
r79 86 93 0.0685365
r80 85 98 0.0685365
r81 85 86 24.7154
r82 52 89 2.16729
r83 47 62 1.16709
r84 47 98 2.12561
r85 43 57 1.16709
r86 43 93 0.5835
r87 40 43 0.0416786
r88 23 57 0.0476429
r89 21 23 0.326018
r90 21 23 0.1167
r91 20 24 0.652036
r92 20 23 6.7686
r93 17 57 0.357321
r94 15 23 0.326018
r95 15 17 0.40845
r96 8 52 1.16709
r97 6 62 0.75
r98 4 24 2.5674
r99 2 17 2.15895
.ends

.subckt PM_G5_XNOR3_N1_VSS 3 6 11 15 18 34 37 44 45 47 54 55 73 78 83 88 93 96
+ 99 108 113 122 124 125 126 131 132 137 145 153 154 155 Vss
c131 155 Vss 3.75522e-19
c132 154 Vss 3.87529e-19
c133 153 Vss 4.4306e-19
c134 137 Vss 0.00333207f
c135 132 Vss 8.38361e-19
c136 131 Vss 0.00578307f
c137 126 Vss 8.35423e-19
c138 125 Vss 0.00509728f
c139 124 Vss 0.0036146f
c140 122 Vss 0.00254978f
c141 113 Vss 0.00381203f
c142 108 Vss 0.0040091f
c143 99 Vss 0.00484046f
c144 96 Vss 0.00348301f
c145 93 Vss 0.00279856f
c146 88 Vss 7.12901e-19
c147 83 Vss 0.00141291f
c148 78 Vss 0.0025656f
c149 73 Vss 0.00249897f
c150 55 Vss 0.0338093f
c151 54 Vss 0.0988897f
c152 47 Vss 7.60188e-20
c153 45 Vss 0.0331638f
c154 44 Vss 0.0974849f
c155 37 Vss 7.50699e-20
c156 35 Vss 0.0349827f
c157 34 Vss 0.1003f
c158 18 Vss 0.00263959f
c159 15 Vss 0.164604f
c160 11 Vss 0.166952f
c161 6 Vss 0.00172036f
c162 3 Vss 0.167004f
r163 143 155 0.494161
r164 143 145 6.71025
r165 139 155 0.128424
r166 138 154 0.494161
r167 137 149 0.652036
r168 137 138 7.46046
r169 133 154 0.128424
r170 131 155 0.494161
r171 131 132 15.8795
r172 127 153 0.0828784
r173 125 154 0.494161
r174 125 126 13.0037
r175 124 132 0.652036
r176 123 153 0.551426
r177 123 124 10.6697
r178 122 153 0.551426
r179 121 126 0.652036
r180 121 122 6.83529
r181 96 145 1.33371
r182 93 96 5.41821
r183 88 113 1.16709
r184 88 149 2.16729
r185 83 108 1.16709
r186 83 139 2.16729
r187 78 133 4.83471
r188 73 99 1.16709
r189 73 127 4.33978
r190 57 113 0.238214
r191 55 57 1.45875
r192 54 58 0.652036
r193 54 57 1.45875
r194 51 55 0.652036
r195 47 108 0.238214
r196 45 47 1.45875
r197 44 48 0.652036
r198 44 47 1.45875
r199 41 45 0.652036
r200 37 99 0.238214
r201 35 37 1.45875
r202 34 38 0.652036
r203 34 37 1.45875
r204 31 35 0.652036
r205 18 93 1.16709
r206 15 58 2.5674
r207 15 51 2.5674
r208 11 48 2.5674
r209 11 41 2.5674
r210 6 78 1.16709
r211 3 38 2.5674
r212 3 31 2.5674
.ends

.subckt PM_G5_XNOR3_N1_CI 2 6 8 34 39 44 79 80 85 91 Vss
c47 91 Vss 2.52123e-19
c48 85 Vss 0.00547442f
c49 80 Vss 3.74154e-19
c50 79 Vss 0.0039666f
c51 44 Vss 0.00209085f
c52 39 Vss 0.00132824f
c53 34 Vss 0.00535743f
c54 8 Vss 0.00276539f
c55 6 Vss 0.00213002f
c56 2 Vss 0.00154503f
r57 86 91 0.494161
r58 85 87 0.652036
r59 85 86 10.3363
r60 81 91 0.128424
r61 79 91 0.494161
r62 79 80 21.8396
r63 75 80 0.652036
r64 44 87 2.16729
r65 39 81 2.16729
r66 34 75 11.3366
r67 8 44 1.16709
r68 6 39 1.16709
r69 2 34 1.16709
.ends

.subckt PM_G5_XNOR3_N1_A 2 4 7 11 21 24 45 49 51 54 56 57 58 62 63 69 74 Vss
c79 74 Vss 0.00491901f
c80 69 Vss 0.00491594f
c81 63 Vss 8.26639e-19
c82 62 Vss 4.20301e-19
c83 58 Vss 0.0011362f
c84 57 Vss 0.00976615f
c85 56 Vss 0.00370619f
c86 51 Vss 0.00520175f
c87 49 Vss 0.135015f
c88 45 Vss 0.126353f
c89 24 Vss 0.2139f
c90 21 Vss 0.0724995f
c91 19 Vss 0.0247918f
c92 7 Vss 1.00425f
c93 4 Vss 0.0850321f
r94 74 77 0.1
r95 66 77 1.16709
r96 63 66 0.833571
r97 60 69 1.16709
r98 60 62 0.513084
r99 57 63 0.0685365
r100 57 58 10.4613
r101 55 58 0.652036
r102 55 56 8.66914
r103 54 62 0.791893
r104 51 56 0.652036
r105 51 54 9.41936
r106 47 49 4.53833
r107 44 74 0.262036
r108 44 45 2.26917
r109 41 44 2.26917
r110 36 49 0.00605528
r111 35 45 0.00605528
r112 32 47 0.00605528
r113 31 41 0.00605528
r114 27 69 0.0952857
r115 25 27 0.326018
r116 25 27 0.1167
r117 24 28 0.652036
r118 24 27 6.7686
r119 21 27 0.3335
r120 19 27 0.326018
r121 19 21 0.2334
r122 11 36 2.5674
r123 11 32 2.5674
r124 7 11 12.837
r125 7 35 2.5674
r126 7 11 12.837
r127 7 31 2.5674
r128 4 28 2.5674
r129 2 21 2.334
.ends

.subckt PM_G5_XNOR3_N1_BI 2 6 8 16 23 32 37 42 51 56 64 65 71 78 83 84 Vss
c70 84 Vss 1.10364e-19
c71 83 Vss 0.00214683f
c72 78 Vss 8.34553e-19
c73 71 Vss 5.02505e-19
c74 65 Vss 4.43116e-19
c75 64 Vss 0.00191151f
c76 56 Vss 0.00250766f
c77 51 Vss 0.00202351f
c78 42 Vss 0.00122467f
c79 37 Vss 4.09629e-19
c80 32 Vss 0.00157267f
c81 23 Vss 7.03109e-20
c82 16 Vss 0.0573997f
c83 8 Vss 0.0573997f
c84 2 Vss 0.00150258f
r85 82 84 0.65228
r86 82 83 3.46076
r87 78 83 0.65228
r88 74 78 2.1006
r89 71 74 2.08393
r90 64 71 0.0685365
r91 64 65 13.2121
r92 60 65 0.652036
r93 42 56 1.16709
r94 42 84 2.1395
r95 37 51 1.16709
r96 37 74 0.0416786
r97 32 60 4.29289
r98 23 56 0.50025
r99 16 51 0.50025
r100 8 23 1.80885
r101 6 16 1.80885
r102 2 32 1.16709
.ends

.subckt PM_G5_XNOR3_N1_AI 2 7 11 31 36 37 46 51 60 69 Vss
c47 69 Vss 2.92061e-19
c48 60 Vss 0.0055297f
c49 51 Vss 0.00389112f
c50 46 Vss 9.98085e-19
c51 37 Vss 0.127837f
c52 36 Vss 5.86204e-20
c53 31 Vss 0.128631f
c54 7 Vss 0.994815f
c55 2 Vss 0.00150258f
r56 65 69 0.652036
r57 60 63 0.1
r58 51 63 1.16709
r59 51 69 13.7539
r60 46 65 2.16729
r61 36 60 0.262036
r62 36 37 2.334
r63 33 36 2.20433
r64 29 31 4.53833
r65 26 37 0.00605528
r66 25 31 0.00605528
r67 22 33 0.00605528
r68 21 29 0.00605528
r69 11 26 2.5674
r70 11 22 2.5674
r71 7 11 12.837
r72 7 25 2.5674
r73 7 11 12.837
r74 7 21 2.5674
r75 2 46 1.16709
.ends

.subckt PM_G5_XNOR3_N1_B 2 4 6 8 16 17 24 28 31 42 45 50 55 60 65 69 76 77 Vss
c63 77 Vss 1.47395e-19
c64 76 Vss 6.32207e-19
c65 69 Vss 0.0035022f
c66 65 Vss 0.00265398f
c67 60 Vss 0.00253939f
c68 55 Vss 0.00274111f
c69 50 Vss 0.00171367f
c70 45 Vss 5.45343e-20
c71 42 Vss 5.46775e-19
c72 31 Vss 0.0573997f
c73 24 Vss 1.2014e-19
c74 20 Vss 0.0247918f
c75 17 Vss 0.0338376f
c76 16 Vss 0.183114f
c77 6 Vss 0.0573997f
c78 4 Vss 0.0714101f
c79 2 Vss 0.0826049f
r80 76 77 0.65228
r81 75 76 3.46076
r82 69 75 0.65228
r83 50 65 1.16709
r84 50 77 2.1395
r85 45 60 1.16709
r86 45 69 2.1006
r87 38 55 1.16709
r88 38 45 10.7364
r89 38 42 0.0364688
r90 36 55 0.0476429
r91 31 65 0.50025
r92 28 60 0.50025
r93 24 55 0.357321
r94 20 36 0.326018
r95 20 24 0.40845
r96 17 36 6.7686
r97 16 36 0.326018
r98 16 36 0.1167
r99 13 17 0.652036
r100 8 31 1.80885
r101 6 28 1.80885
r102 4 24 2.15895
r103 2 13 2.5674
.ends

.subckt PM_G5_XNOR3_N1_Z 2 4 30 33 Vss
c31 30 Vss 0.00315811f
c32 4 Vss 0.00153036f
c33 2 Vss 0.00166246f
r34 33 35 4.20954
r35 30 33 4.95975
r36 4 35 1.16709
r37 2 30 1.16709
.ends

.subckt G5_XNOR3_N1  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI10.X0 N_CI_XI10.X0_D N_VSS_XI10.X0_PGD N_C_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW4
XI9.X0 N_CI_XI10.X0_D N_VDD_XI9.X0_PGD N_C_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI5.X0 N_BI_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI6.X0 N_BI_XI5.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW4
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW4
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_B_XI2.X0_CG N_AI_XI2.X0_PGD N_C_XI2.X0_S
+ TIGFET_HPNW4
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_BI_XI4.X0_CG N_AI_XI4.X0_PGD N_CI_XI4.X0_S
+ TIGFET_HPNW4
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_BI_XI3.X0_CG N_A_XI3.X0_PGD N_C_XI3.X0_S
+ TIGFET_HPNW4
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_B_XI1.X0_CG N_A_XI1.X0_PGD N_CI_XI1.X0_S
+ TIGFET_HPNW4
*
x_PM_G5_XNOR3_N1_VDD N_VDD_XI10.X0_S N_VDD_XI9.X0_PGD N_VDD_XI5.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI6.X0_S N_VDD_XI7.X0_PGD N_VDD_c_120_p N_VDD_c_18_p
+ N_VDD_c_23_p N_VDD_c_4_p N_VDD_c_110_p N_VDD_c_19_p N_VDD_c_6_p N_VDD_c_25_p
+ N_VDD_c_5_p N_VDD_c_64_p N_VDD_c_27_p N_VDD_c_28_p N_VDD_c_29_p N_VDD_c_35_p
+ N_VDD_c_32_p N_VDD_c_20_p N_VDD_c_11_p N_VDD_c_24_p N_VDD_c_37_p N_VDD_c_12_p
+ N_VDD_c_60_p VDD N_VDD_c_68_p N_VDD_c_72_p N_VDD_c_2_p N_VDD_c_42_p
+ N_VDD_c_38_p Vss PM_G5_XNOR3_N1_VDD
x_PM_G5_XNOR3_N1_C N_C_XI10.X0_CG N_C_XI9.X0_CG N_C_XI2.X0_S N_C_XI3.X0_S
+ N_C_c_143_p N_C_c_125_n N_C_c_136_p C N_C_c_138_p N_C_c_158_p N_C_c_178_p
+ N_C_c_130_n N_C_c_132_n N_C_c_133_n N_C_c_156_p N_C_c_139_p N_C_c_161_p Vss
+ PM_G5_XNOR3_N1_C
x_PM_G5_XNOR3_N1_VSS N_VSS_XI10.X0_PGD N_VSS_XI9.X0_S N_VSS_XI8.X0_PGD
+ N_VSS_XI6.X0_PGD N_VSS_XI7.X0_S N_VSS_c_188_n N_VSS_c_247_n N_VSS_c_189_n
+ N_VSS_c_191_n N_VSS_c_287_p N_VSS_c_192_n N_VSS_c_193_n N_VSS_c_195_n
+ N_VSS_c_201_n N_VSS_c_205_n N_VSS_c_209_n N_VSS_c_213_n N_VSS_c_216_n
+ N_VSS_c_217_n N_VSS_c_220_n N_VSS_c_224_n N_VSS_c_228_n N_VSS_c_231_n
+ N_VSS_c_233_n N_VSS_c_234_n N_VSS_c_235_n N_VSS_c_239_n N_VSS_c_240_n VSS
+ N_VSS_c_243_n N_VSS_c_244_n N_VSS_c_245_n Vss PM_G5_XNOR3_N1_VSS
x_PM_G5_XNOR3_N1_CI N_CI_XI10.X0_D N_CI_XI4.X0_S N_CI_XI1.X0_S N_CI_c_316_n
+ N_CI_c_334_n N_CI_c_356_p N_CI_c_320_n N_CI_c_338_n N_CI_c_324_n N_CI_c_349_p
+ Vss PM_G5_XNOR3_N1_CI
x_PM_G5_XNOR3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI3.X0_PGD N_A_XI1.X0_PGD
+ N_A_c_387_n N_A_c_362_n N_A_c_415_p N_A_c_417_p N_A_c_363_n A N_A_c_370_n
+ N_A_c_381_n N_A_c_371_n N_A_c_372_n N_A_c_386_n N_A_c_374_n N_A_c_399_p Vss
+ PM_G5_XNOR3_N1_A
x_PM_G5_XNOR3_N1_BI N_BI_XI5.X0_D N_BI_XI4.X0_CG N_BI_XI3.X0_CG N_BI_c_478_p
+ N_BI_c_465_n N_BI_c_443_n N_BI_c_468_n N_BI_c_459_n N_BI_c_471_n N_BI_c_472_n
+ N_BI_c_447_n N_BI_c_457_n N_BI_c_477_n N_BI_c_450_n N_BI_c_503_p N_BI_c_451_n
+ Vss PM_G5_XNOR3_N1_BI
x_PM_G5_XNOR3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_523_n
+ N_AI_c_546_n N_AI_c_513_n N_AI_c_514_n N_AI_c_517_n N_AI_c_528_n N_AI_c_518_n
+ Vss PM_G5_XNOR3_N1_AI
x_PM_G5_XNOR3_N1_B N_B_XI5.X0_CG N_B_XI6.X0_CG N_B_XI2.X0_CG N_B_XI1.X0_CG
+ N_B_c_559_n N_B_c_561_n N_B_c_571_n N_B_c_580_n N_B_c_581_n B N_B_c_584_n
+ N_B_c_575_n N_B_c_562_n N_B_c_589_n N_B_c_590_n N_B_c_563_n N_B_c_607_n
+ N_B_c_576_n Vss PM_G5_XNOR3_N1_B
x_PM_G5_XNOR3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_624_n Z Vss PM_G5_XNOR3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_C_XI9.X0_CG 9.58934e-19
cc_2 N_VDD_c_2_p N_C_XI9.X0_CG 8.03148e-19
cc_3 N_VDD_XI9.X0_PGD N_C_c_125_n 4.16623e-19
cc_4 N_VDD_c_4_p N_C_c_125_n 9.58934e-19
cc_5 N_VDD_c_5_p N_C_c_125_n 0.00125128f
cc_6 N_VDD_c_6_p C 3.00172e-19
cc_7 N_VDD_c_5_p C 0.00118142f
cc_8 N_VDD_c_6_p N_C_c_130_n 4.71537e-19
cc_9 N_VDD_c_5_p N_C_c_130_n 2.74773e-19
cc_10 N_VDD_XI6.X0_S N_C_c_132_n 3.43419e-19
cc_11 N_VDD_c_11_p N_C_c_133_n 5.30636e-19
cc_12 N_VDD_c_12_p N_C_c_133_n 7.99481e-19
cc_13 N_VDD_XI9.X0_PGD N_VSS_XI10.X0_PGD 0.00173038f
cc_14 N_VDD_XI5.X0_PGD N_VSS_XI8.X0_PGD 2.27468e-19
cc_15 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172039f
cc_16 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017188f
cc_17 N_VDD_XI7.X0_PGD N_VSS_XI6.X0_PGD 2.1536e-19
cc_18 N_VDD_c_18_p N_VSS_c_188_n 0.00173038f
cc_19 N_VDD_c_19_p N_VSS_c_189_n 0.00172039f
cc_20 N_VDD_c_20_p N_VSS_c_189_n 2.46461e-19
cc_21 N_VDD_c_20_p N_VSS_c_191_n 3.60588e-19
cc_22 N_VDD_c_12_p N_VSS_c_192_n 2.35445e-19
cc_23 N_VDD_c_23_p N_VSS_c_193_n 0.0017188f
cc_24 N_VDD_c_24_p N_VSS_c_193_n 2.74208e-19
cc_25 N_VDD_c_25_p N_VSS_c_195_n 4.32468e-19
cc_26 N_VDD_c_5_p N_VSS_c_195_n 4.60511e-19
cc_27 N_VDD_c_27_p N_VSS_c_195_n 0.00130521f
cc_28 N_VDD_c_28_p N_VSS_c_195_n 4.50568e-19
cc_29 N_VDD_c_29_p N_VSS_c_195_n 3.98949e-19
cc_30 N_VDD_c_2_p N_VSS_c_195_n 3.48267e-19
cc_31 N_VDD_c_5_p N_VSS_c_201_n 5.01863e-19
cc_32 N_VDD_c_32_p N_VSS_c_201_n 2.14355e-19
cc_33 N_VDD_c_11_p N_VSS_c_201_n 7.9087e-19
cc_34 N_VDD_c_12_p N_VSS_c_201_n 3.30117e-19
cc_35 N_VDD_c_35_p N_VSS_c_205_n 6.99368e-19
cc_36 N_VDD_c_20_p N_VSS_c_205_n 0.00161703f
cc_37 N_VDD_c_37_p N_VSS_c_205_n 8.32098e-19
cc_38 N_VDD_c_38_p N_VSS_c_205_n 3.48267e-19
cc_39 N_VDD_c_11_p N_VSS_c_209_n 6.79271e-19
cc_40 N_VDD_c_24_p N_VSS_c_209_n 0.00161703f
cc_41 N_VDD_c_12_p N_VSS_c_209_n 0.00241473f
cc_42 N_VDD_c_42_p N_VSS_c_209_n 3.48267e-19
cc_43 N_VDD_XI7.X0_PGD N_VSS_c_213_n 3.41313e-19
cc_44 N_VDD_c_37_p N_VSS_c_213_n 0.00506009f
cc_45 N_VDD_c_38_p N_VSS_c_213_n 9.58524e-19
cc_46 N_VDD_c_20_p N_VSS_c_216_n 0.00415364f
cc_47 N_VDD_c_25_p N_VSS_c_217_n 4.41003e-19
cc_48 N_VDD_c_29_p N_VSS_c_217_n 3.89161e-19
cc_49 N_VDD_c_2_p N_VSS_c_217_n 7.99831e-19
cc_50 N_VDD_c_35_p N_VSS_c_220_n 3.48267e-19
cc_51 N_VDD_c_20_p N_VSS_c_220_n 2.03837e-19
cc_52 N_VDD_c_37_p N_VSS_c_220_n 3.99794e-19
cc_53 N_VDD_c_38_p N_VSS_c_220_n 8.03027e-19
cc_54 N_VDD_c_11_p N_VSS_c_224_n 3.82294e-19
cc_55 N_VDD_c_24_p N_VSS_c_224_n 2.03837e-19
cc_56 N_VDD_c_12_p N_VSS_c_224_n 9.55109e-19
cc_57 N_VDD_c_42_p N_VSS_c_224_n 8.01441e-19
cc_58 N_VDD_c_6_p N_VSS_c_228_n 0.00301593f
cc_59 N_VDD_c_25_p N_VSS_c_228_n 7.60301e-19
cc_60 N_VDD_c_60_p N_VSS_c_228_n 0.0010705f
cc_61 N_VDD_c_25_p N_VSS_c_231_n 0.00803422f
cc_62 N_VDD_c_29_p N_VSS_c_231_n 8.94414e-19
cc_63 N_VDD_c_5_p N_VSS_c_233_n 0.00969041f
cc_64 N_VDD_c_64_p N_VSS_c_234_n 0.00107143f
cc_65 N_VDD_c_28_p N_VSS_c_235_n 0.00807788f
cc_66 N_VDD_c_32_p N_VSS_c_235_n 7.22996e-19
cc_67 N_VDD_c_20_p N_VSS_c_235_n 0.00374557f
cc_68 N_VDD_c_68_p N_VSS_c_235_n 0.00137227f
cc_69 N_VDD_c_25_p N_VSS_c_239_n 0.00107355f
cc_70 N_VDD_c_5_p N_VSS_c_240_n 0.00142851f
cc_71 N_VDD_c_24_p N_VSS_c_240_n 0.00577339f
cc_72 N_VDD_c_72_p N_VSS_c_240_n 0.00106333f
cc_73 N_VDD_c_25_p N_VSS_c_243_n 0.00112682f
cc_74 N_VDD_c_5_p N_VSS_c_244_n 0.00104966f
cc_75 N_VDD_c_20_p N_VSS_c_245_n 7.74609e-19
cc_76 N_VDD_XI10.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_77 N_VDD_c_27_p N_CI_XI10.X0_D 3.72199e-19
cc_78 N_VDD_XI10.X0_S N_CI_c_316_n 3.48267e-19
cc_79 N_VDD_c_5_p N_CI_c_316_n 5.01863e-19
cc_80 N_VDD_c_27_p N_CI_c_316_n 5.226e-19
cc_81 N_VDD_c_29_p N_CI_c_316_n 0.00213742f
cc_82 N_VDD_c_35_p N_CI_c_320_n 7.47076e-19
cc_83 N_VDD_c_32_p N_CI_c_320_n 4.06004e-19
cc_84 N_VDD_c_38_p N_A_XI7.X0_CG 9.92565e-19
cc_85 N_VDD_XI7.X0_PGD N_A_c_362_n 3.90792e-19
cc_86 N_VDD_XI6.X0_S N_A_c_363_n 2.96819e-19
cc_87 N_VDD_XI7.X0_PGD N_A_c_363_n 5.17967e-19
cc_88 N_VDD_c_20_p N_A_c_363_n 4.32724e-19
cc_89 N_VDD_c_24_p N_A_c_363_n 4.10602e-19
cc_90 N_VDD_c_37_p N_A_c_363_n 4.1682e-19
cc_91 N_VDD_c_12_p N_A_c_363_n 3.91173e-19
cc_92 N_VDD_c_38_p N_A_c_363_n 5.53168e-19
cc_93 N_VDD_XI6.X0_S N_A_c_370_n 9.18655e-19
cc_94 N_VDD_c_12_p N_A_c_371_n 0.00608947f
cc_95 N_VDD_c_29_p N_A_c_372_n 8.16868e-19
cc_96 N_VDD_c_11_p N_A_c_372_n 2.36389e-19
cc_97 N_VDD_c_29_p N_A_c_374_n 6.33536e-19
cc_98 N_VDD_c_42_p N_A_c_374_n 5.39283e-19
cc_99 N_VDD_XI6.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_100 N_VDD_c_24_p N_BI_XI5.X0_D 3.7884e-19
cc_101 N_VDD_c_12_p N_BI_XI5.X0_D 3.48267e-19
cc_102 N_VDD_XI6.X0_S N_BI_c_443_n 3.48267e-19
cc_103 N_VDD_c_29_p N_BI_c_443_n 8.52765e-19
cc_104 N_VDD_c_24_p N_BI_c_443_n 4.58491e-19
cc_105 N_VDD_c_12_p N_BI_c_443_n 7.03408e-19
cc_106 N_VDD_c_24_p N_BI_c_447_n 2.4324e-19
cc_107 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_108 N_VDD_c_32_p N_AI_XI8.X0_D 3.73302e-19
cc_109 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.86706e-19
cc_110 N_VDD_c_110_p N_AI_c_513_n 2.86706e-19
cc_111 N_VDD_XI8.X0_S N_AI_c_514_n 3.48267e-19
cc_112 N_VDD_c_32_p N_AI_c_514_n 5.23123e-19
cc_113 N_VDD_c_20_p N_AI_c_514_n 5.01863e-19
cc_114 N_VDD_c_37_p N_AI_c_517_n 0.00111556f
cc_115 N_VDD_c_20_p N_AI_c_518_n 2.2965e-19
cc_116 N_VDD_XI9.X0_PGD N_B_XI5.X0_CG 9.5906e-19
cc_117 N_VDD_c_42_p N_B_XI5.X0_CG 9.74645e-19
cc_118 N_VDD_XI5.X0_PGD N_B_c_559_n 3.9688e-19
cc_119 N_VDD_XI7.X0_PGD N_B_c_559_n 2.07132e-19
cc_120 N_VDD_c_120_p N_B_c_561_n 9.5906e-19
cc_121 N_VDD_c_38_p N_B_c_562_n 2.92921e-19
cc_122 N_VDD_c_12_p N_B_c_563_n 5.34599e-19
cc_123 N_C_c_125_n N_VSS_XI10.X0_PGD 4.16623e-19
cc_124 N_C_c_136_p N_VSS_c_247_n 9.33417e-19
cc_125 C N_VSS_c_195_n 6.06998e-19
cc_126 N_C_c_138_p N_VSS_c_195_n 4.82229e-19
cc_127 N_C_c_139_p N_VSS_c_195_n 2.78014e-19
cc_128 N_C_c_138_p N_VSS_c_201_n 2.30642e-19
cc_129 N_C_c_133_n N_VSS_c_201_n 0.00197293f
cc_130 N_C_c_133_n N_VSS_c_209_n 0.00165406f
cc_131 N_C_c_143_p N_VSS_c_217_n 0.0041205f
cc_132 N_C_c_136_p N_VSS_c_217_n 7.00195e-19
cc_133 C N_VSS_c_217_n 4.56568e-19
cc_134 N_C_c_130_n N_VSS_c_217_n 6.1245e-19
cc_135 C N_VSS_c_228_n 2.17246e-19
cc_136 N_C_c_138_p N_VSS_c_228_n 4.01014e-19
cc_137 N_C_c_139_p N_VSS_c_228_n 4.34874e-19
cc_138 C N_VSS_c_233_n 2.70819e-19
cc_139 N_C_c_138_p N_VSS_c_233_n 9.65301e-19
cc_140 N_C_c_139_p N_VSS_c_233_n 0.00282977f
cc_141 N_C_c_133_n N_VSS_c_240_n 0.00175198f
cc_142 N_C_c_133_n N_CI_c_316_n 0.00136327f
cc_143 N_C_c_133_n N_CI_c_320_n 0.00242327f
cc_144 N_C_c_156_p N_CI_c_324_n 4.1018e-19
cc_145 N_C_c_133_n N_A_c_363_n 2.5075e-19
cc_146 N_C_c_158_p N_A_c_370_n 0.00148519f
cc_147 N_C_c_132_n N_A_c_370_n 8.20481e-19
cc_148 N_C_c_133_n N_A_c_370_n 2.96346e-19
cc_149 N_C_c_161_p N_A_c_370_n 2.4205e-19
cc_150 N_C_c_158_p N_A_c_381_n 0.00189731f
cc_151 N_C_c_132_n N_A_c_381_n 9.00742e-19
cc_152 N_C_c_133_n N_A_c_381_n 3.9734e-19
cc_153 N_C_c_156_p N_A_c_381_n 0.00207353f
cc_154 N_C_c_161_p N_A_c_381_n 6.32429e-19
cc_155 N_C_c_156_p N_A_c_386_n 5.4333e-19
cc_156 N_C_c_133_n N_BI_c_443_n 2.41407e-19
cc_157 N_C_c_133_n N_BI_c_447_n 4.13621e-19
cc_158 N_C_c_156_p N_BI_c_450_n 6.74177e-19
cc_159 N_C_c_156_p N_BI_c_451_n 0.00240592f
cc_160 N_C_c_158_p N_B_c_563_n 0.00168372f
cc_161 N_C_c_133_n N_B_c_563_n 0.0027048f
cc_162 N_C_c_156_p N_B_c_563_n 0.00182275f
cc_163 N_C_c_161_p N_B_c_563_n 2.1095e-19
cc_164 N_C_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_165 N_C_c_158_p N_Z_XI2.X0_D 3.48267e-19
cc_166 N_C_c_178_p N_Z_XI2.X0_D 3.48267e-19
cc_167 N_C_c_132_n N_Z_XI2.X0_D 3.43419e-19
cc_168 N_C_XI3.X0_S N_Z_c_624_n 3.48267e-19
cc_169 N_C_c_158_p N_Z_c_624_n 3.41702e-19
cc_170 N_C_c_178_p N_Z_c_624_n 5.7093e-19
cc_171 N_VSS_XI9.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_172 N_VSS_c_201_n N_CI_XI10.X0_D 3.48267e-19
cc_173 N_VSS_XI7.X0_S N_CI_XI4.X0_S 3.43419e-19
cc_174 N_VSS_c_213_n N_CI_XI4.X0_S 3.48267e-19
cc_175 N_VSS_XI9.X0_S N_CI_c_316_n 3.48267e-19
cc_176 N_VSS_c_195_n N_CI_c_316_n 5.78167e-19
cc_177 N_VSS_c_201_n N_CI_c_316_n 0.00107566f
cc_178 N_VSS_c_231_n N_CI_c_316_n 0.0020072f
cc_179 N_VSS_c_233_n N_CI_c_316_n 3.32126e-19
cc_180 N_VSS_XI7.X0_S N_CI_c_334_n 3.48267e-19
cc_181 N_VSS_c_213_n N_CI_c_334_n 9.13167e-19
cc_182 N_VSS_c_205_n N_CI_c_320_n 0.00134034f
cc_183 N_VSS_c_216_n N_CI_c_320_n 0.00393483f
cc_184 N_VSS_c_235_n N_CI_c_338_n 0.00292666f
cc_185 N_VSS_c_220_n N_A_c_387_n 0.00236445f
cc_186 N_VSS_XI8.X0_PGD N_A_c_362_n 3.86211e-19
cc_187 N_VSS_XI7.X0_S N_A_c_363_n 9.18655e-19
cc_188 N_VSS_c_213_n N_A_c_363_n 0.00149545f
cc_189 N_VSS_c_216_n N_A_c_363_n 2.12774e-19
cc_190 N_VSS_c_240_n N_A_c_363_n 2.27118e-19
cc_191 N_VSS_c_205_n N_A_c_372_n 4.58305e-19
cc_192 N_VSS_c_220_n N_A_c_372_n 4.30193e-19
cc_193 N_VSS_c_287_p N_A_c_374_n 8.53264e-19
cc_194 N_VSS_c_205_n N_A_c_374_n 4.26083e-19
cc_195 N_VSS_c_220_n N_A_c_374_n 7.20776e-19
cc_196 N_VSS_XI9.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_197 N_VSS_c_201_n N_BI_XI5.X0_D 3.48267e-19
cc_198 N_VSS_XI9.X0_S N_BI_c_443_n 3.48267e-19
cc_199 N_VSS_c_201_n N_BI_c_443_n 0.00102079f
cc_200 N_VSS_c_240_n N_BI_c_443_n 3.31365e-19
cc_201 N_VSS_c_216_n N_BI_c_457_n 2.90278e-19
cc_202 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_203 N_VSS_c_213_n N_AI_XI8.X0_D 3.48267e-19
cc_204 N_VSS_XI6.X0_PGD N_AI_XI2.X0_PGD 2.84687e-19
cc_205 N_VSS_c_213_n N_AI_XI2.X0_PGD 2.04949e-19
cc_206 N_VSS_c_192_n N_AI_c_523_n 2.84687e-19
cc_207 N_VSS_XI7.X0_S N_AI_c_514_n 3.48267e-19
cc_208 N_VSS_c_205_n N_AI_c_514_n 0.00163244f
cc_209 N_VSS_c_213_n N_AI_c_514_n 0.00129029f
cc_210 N_VSS_c_213_n N_AI_c_517_n 0.00168777f
cc_211 N_VSS_c_213_n N_AI_c_528_n 2.82216e-19
cc_212 N_VSS_c_216_n N_AI_c_518_n 0.00857137f
cc_213 N_VSS_c_224_n N_B_XI6.X0_CG 0.00272012f
cc_214 N_VSS_XI8.X0_PGD N_B_c_559_n 2.07132e-19
cc_215 N_VSS_XI6.X0_PGD N_B_c_559_n 3.923e-19
cc_216 N_VSS_c_224_n N_B_c_571_n 0.00138168f
cc_217 N_VSS_c_209_n B 5.92764e-19
cc_218 N_VSS_c_224_n N_B_c_562_n 6.1245e-19
cc_219 N_VSS_c_209_n N_B_c_563_n 6.44904e-19
cc_220 N_CI_c_316_n N_BI_c_443_n 0.00104494f
cc_221 N_CI_c_324_n N_BI_c_459_n 6.86101e-19
cc_222 N_CI_c_334_n N_BI_c_447_n 8.7e-19
cc_223 N_CI_c_320_n N_BI_c_447_n 9.27611e-19
cc_224 N_CI_c_324_n N_BI_c_450_n 0.00228179f
cc_225 N_CI_c_316_n N_AI_c_514_n 5.24832e-19
cc_226 N_CI_c_334_n N_AI_c_514_n 5.10362e-19
cc_227 N_CI_c_334_n N_AI_c_517_n 0.00202744f
cc_228 N_CI_c_320_n N_AI_c_517_n 0.00654866f
cc_229 N_CI_c_324_n N_AI_c_517_n 0.00288502f
cc_230 N_CI_c_349_p N_AI_c_517_n 8.49574e-19
cc_231 N_CI_c_320_n N_AI_c_518_n 9.37419e-19
cc_232 N_CI_c_324_n N_B_c_575_n 0.00103435f
cc_233 N_CI_c_324_n N_B_c_576_n 2.42418e-19
cc_234 N_CI_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_235 N_CI_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_236 N_CI_c_334_n N_Z_XI4.X0_D 3.48267e-19
cc_237 N_CI_c_356_p N_Z_XI4.X0_D 3.48267e-19
cc_238 N_CI_XI4.X0_S N_Z_c_624_n 3.48267e-19
cc_239 N_CI_XI1.X0_S N_Z_c_624_n 3.48267e-19
cc_240 N_CI_c_334_n N_Z_c_624_n 5.68744e-19
cc_241 N_CI_c_356_p N_Z_c_624_n 5.68744e-19
cc_242 N_A_XI3.X0_PGD N_BI_XI3.X0_CG 8.79767e-19
cc_243 N_A_c_399_p N_BI_XI3.X0_CG 0.00237738f
cc_244 N_A_c_399_p N_BI_c_465_n 0.00117691f
cc_245 N_A_c_363_n N_BI_c_443_n 4.0484e-19
cc_246 N_A_c_370_n N_BI_c_443_n 6.63236e-19
cc_247 N_A_c_363_n N_BI_c_468_n 2.37396e-19
cc_248 N_A_c_386_n N_BI_c_459_n 7.92141e-19
cc_249 N_A_c_399_p N_BI_c_459_n 4.87897e-19
cc_250 N_A_c_363_n N_BI_c_471_n 3.8563e-19
cc_251 N_A_XI3.X0_PGD N_BI_c_472_n 0.00133285f
cc_252 N_A_c_386_n N_BI_c_472_n 4.79282e-19
cc_253 N_A_c_399_p N_BI_c_472_n 0.00152548f
cc_254 N_A_c_370_n N_BI_c_447_n 0.00181644f
cc_255 N_A_c_363_n N_BI_c_457_n 0.00247154f
cc_256 N_A_c_370_n N_BI_c_477_n 2.27623e-19
cc_257 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174824f
cc_258 N_A_c_370_n N_AI_XI2.X0_PGD 8.597e-19
cc_259 N_A_c_415_p N_AI_c_523_n 0.00199346f
cc_260 N_A_c_381_n N_AI_c_523_n 0.00123218f
cc_261 N_A_c_417_p N_AI_c_513_n 0.00202303f
cc_262 N_A_c_363_n N_AI_c_514_n 0.00165136f
cc_263 N_A_c_363_n N_AI_c_517_n 0.00184834f
cc_264 N_A_c_362_n N_B_c_559_n 0.00360254f
cc_265 N_A_c_363_n N_B_c_559_n 5.41329e-19
cc_266 N_A_c_374_n N_B_c_561_n 4.14098e-19
cc_267 N_A_c_381_n N_B_c_580_n 2.74862e-19
cc_268 N_A_XI3.X0_PGD N_B_c_581_n 8.79767e-19
cc_269 N_A_c_363_n B 6.972e-19
cc_270 N_A_c_370_n B 3.89684e-19
cc_271 N_A_c_370_n N_B_c_584_n 3.55503e-19
cc_272 N_A_c_381_n N_B_c_584_n 4.94081e-19
cc_273 N_A_c_381_n N_B_c_575_n 3.26384e-19
cc_274 N_A_c_362_n N_B_c_562_n 2.86506e-19
cc_275 N_A_c_370_n N_B_c_562_n 6.34732e-19
cc_276 N_A_c_370_n N_B_c_589_n 3.37713e-19
cc_277 N_A_XI3.X0_PGD N_B_c_590_n 0.00133285f
cc_278 N_A_c_370_n N_B_c_563_n 0.00206097f
cc_279 N_A_c_381_n N_B_c_563_n 0.00238641f
cc_280 N_A_c_381_n N_Z_XI2.X0_D 6.94686e-19
cc_281 N_A_XI3.X0_PGD N_Z_c_624_n 6.45939e-19
cc_282 N_A_c_370_n N_Z_c_624_n 0.00131646f
cc_283 N_A_c_381_n N_Z_c_624_n 0.00121415f
cc_284 N_BI_c_478_p N_AI_XI2.X0_PGD 8.79767e-19
cc_285 N_BI_c_471_n N_AI_XI2.X0_PGD 0.00133285f
cc_286 N_BI_c_471_n N_AI_c_546_n 6.37981e-19
cc_287 N_BI_c_457_n N_AI_c_514_n 8.05284e-19
cc_288 N_BI_c_468_n N_AI_c_517_n 4.93364e-19
cc_289 N_BI_c_447_n N_AI_c_517_n 0.00402897f
cc_290 N_BI_c_477_n N_AI_c_517_n 4.42808e-19
cc_291 N_BI_c_478_p N_AI_c_528_n 0.00234569f
cc_292 N_BI_c_468_n N_AI_c_528_n 4.6759e-19
cc_293 N_BI_c_471_n N_AI_c_528_n 0.00166302f
cc_294 N_BI_c_443_n B 4.30856e-19
cc_295 N_BI_c_447_n B 3.14738e-19
cc_296 N_BI_c_468_n N_B_c_584_n 5.92939e-19
cc_297 N_BI_c_477_n N_B_c_584_n 3.24098e-19
cc_298 N_BI_c_459_n N_B_c_575_n 0.0018551f
cc_299 N_BI_c_471_n N_B_c_589_n 0.00266367f
cc_300 N_BI_c_472_n N_B_c_589_n 6.17967e-19
cc_301 N_BI_c_471_n N_B_c_590_n 7.16621e-19
cc_302 N_BI_c_472_n N_B_c_590_n 0.00243799f
cc_303 N_BI_c_443_n N_B_c_563_n 0.00165434f
cc_304 N_BI_c_459_n N_B_c_563_n 0.00159414f
cc_305 N_BI_c_447_n N_B_c_563_n 0.0157983f
cc_306 N_BI_c_450_n N_B_c_563_n 6.88876e-19
cc_307 N_BI_c_451_n N_B_c_563_n 8.27361e-19
cc_308 N_BI_c_477_n N_B_c_607_n 0.00346365f
cc_309 N_BI_c_503_p N_B_c_607_n 0.00194674f
cc_310 N_BI_c_468_n N_B_c_576_n 3.02576e-19
cc_311 N_BI_c_450_n N_B_c_576_n 8.19447e-19
cc_312 N_BI_c_468_n N_Z_c_624_n 0.00155391f
cc_313 N_BI_c_459_n N_Z_c_624_n 0.00136914f
cc_314 N_BI_c_472_n N_Z_c_624_n 8.66889e-19
cc_315 N_BI_c_477_n N_Z_c_624_n 4.81308e-19
cc_316 N_AI_XI2.X0_PGD N_B_XI2.X0_CG 8.63152e-19
cc_317 N_AI_XI2.X0_PGD N_B_c_589_n 0.00133285f
cc_318 N_AI_XI2.X0_PGD N_Z_c_624_n 3.30612e-19
cc_319 N_B_c_584_n N_Z_c_624_n 0.00130267f
cc_320 N_B_c_575_n N_Z_c_624_n 0.00130267f
cc_321 N_B_c_589_n N_Z_c_624_n 8.66889e-19
cc_322 N_B_c_590_n N_Z_c_624_n 8.66889e-19
cc_323 N_B_c_563_n N_Z_c_624_n 0.00103251f
cc_324 N_B_c_607_n N_Z_c_624_n 0.00216955f
cc_325 N_B_c_576_n N_Z_c_624_n 9.92382e-19
*
.ends
*
*
.subckt XNOR3_HPNW4 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XNOR3_N1
.ends
*
* File: G4_XOR2_N1.pex.netlist
* Created: Fri Mar 18 15:34:38 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XOR2_N1_VSS 2 5 9 12 16 32 33 35 42 43 66 71 76 81 86 95 100 113
+ 115 116 117 122 123 128 138 140 145 146 147 150 Vss
c105 148 Vss 6.13404e-19
c106 147 Vss 3.75522e-19
c107 146 Vss 4.28045e-19
c108 145 Vss 0.0035844f
c109 140 Vss 0.00192576f
c110 138 Vss 0.00847727f
c111 128 Vss 0.00326939f
c112 123 Vss 8.39752e-19
c113 122 Vss 0.00163882f
c114 117 Vss 8.17785e-19
c115 116 Vss 0.00399757f
c116 115 Vss 0.00448448f
c117 113 Vss 0.00145652f
c118 100 Vss 0.00421853f
c119 95 Vss 0.00425358f
c120 86 Vss 1.76201e-20
c121 81 Vss 0.00164759f
c122 76 Vss 7.42069e-19
c123 71 Vss 9.70701e-19
c124 66 Vss 0.0014444f
c125 43 Vss 0.033325f
c126 42 Vss 0.0990681f
c127 35 Vss 7.82991e-20
c128 33 Vss 0.0341879f
c129 32 Vss 0.0981149f
c130 16 Vss 0.00276316f
c131 12 Vss 0.00263275f
c132 9 Vss 0.165244f
c133 5 Vss 0.166856f
c134 2 Vss 0.00267051f
r135 145 150 0.326018
r136 144 145 4.16786
r137 140 144 0.655813
r138 139 148 0.494161
r139 138 150 0.326018
r140 138 139 13.0037
r141 134 148 0.128424
r142 129 147 0.494161
r143 128 148 0.494161
r144 128 129 7.46046
r145 124 147 0.128424
r146 122 147 0.494161
r147 122 123 4.37625
r148 118 146 0.0828784
r149 116 130 0.652036
r150 116 117 10.1279
r151 115 123 0.652036
r152 114 146 0.551426
r153 114 115 12.4619
r154 113 146 0.551426
r155 112 117 0.652036
r156 112 113 4.16786
r157 86 140 1.82344
r158 81 134 4.83471
r159 76 100 1.16709
r160 76 130 2.16729
r161 71 95 1.16709
r162 71 124 2.16729
r163 66 118 1.82344
r164 45 100 0.238214
r165 43 45 1.45875
r166 42 46 0.652036
r167 42 45 1.45875
r168 39 43 0.652036
r169 35 95 0.238214
r170 33 35 1.45875
r171 32 36 0.652036
r172 32 35 1.45875
r173 29 33 0.652036
r174 16 86 1.16709
r175 12 81 1.16709
r176 9 46 2.5674
r177 9 39 2.5674
r178 5 36 2.5674
r179 5 29 2.5674
r180 2 66 1.16709
.ends

.subckt PM_G4_XOR2_N1_VDD 3 6 8 11 16 32 42 43 66 68 69 70 73 75 76 79 81 85 89
+ 91 93 98 99 100 103 109 114 Vss
c106 114 Vss 0.00542312f
c107 109 Vss 0.00583104f
c108 101 Vss 8.76285e-19
c109 100 Vss 2.39889e-19
c110 99 Vss 3.56526e-19
c111 98 Vss 0.00433275f
c112 93 Vss 0.00130328f
c113 91 Vss 0.0132502f
c114 89 Vss 0.0018632f
c115 85 Vss 7.3942e-19
c116 81 Vss 0.00447795f
c117 79 Vss 0.00129126f
c118 76 Vss 8.63329e-19
c119 75 Vss 0.00575889f
c120 73 Vss 0.00159649f
c121 70 Vss 8.67402e-19
c122 69 Vss 0.00219856f
c123 68 Vss 0.00201914f
c124 66 Vss 0.0065263f
c125 43 Vss 0.0341287f
c126 42 Vss 0.099962f
c127 33 Vss 0.0348624f
c128 32 Vss 0.0999592f
c129 16 Vss 0.00189547f
c130 11 Vss 0.165401f
c131 8 Vss 0.00162509f
c132 6 Vss 0.00218552f
c133 3 Vss 0.165774f
r134 98 103 0.349767
r135 97 98 4.16786
r136 93 103 0.306046
r137 93 95 1.82344
r138 92 101 0.494161
r139 91 97 0.652036
r140 91 92 13.0037
r141 87 101 0.128424
r142 87 89 4.83471
r143 85 114 1.16709
r144 83 85 2.16729
r145 82 100 0.494161
r146 81 101 0.494161
r147 81 82 7.46046
r148 79 109 1.16709
r149 77 100 0.128424
r150 77 79 2.16729
r151 75 83 0.652036
r152 75 76 10.1279
r153 71 99 0.0828784
r154 71 73 1.82344
r155 69 100 0.494161
r156 69 70 4.37625
r157 68 76 0.652036
r158 67 99 0.551426
r159 67 68 4.16786
r160 66 99 0.551426
r161 65 70 0.652036
r162 65 66 12.4619
r163 45 114 0.238214
r164 43 45 1.45875
r165 42 46 0.652036
r166 42 45 1.45875
r167 39 43 0.652036
r168 35 109 0.238214
r169 33 35 1.45875
r170 32 36 0.652036
r171 32 35 1.45875
r172 29 33 0.652036
r173 16 95 1.16709
r174 11 46 2.5674
r175 11 39 2.5674
r176 8 89 1.16709
r177 6 73 1.02121
r178 3 36 2.5674
r179 3 29 2.5674
.ends

.subckt PM_G4_XOR2_N1_A 2 4 7 10 18 21 24 28 39 48 54 57 62 67 72 77 85 Vss
c59 85 Vss 4.11933e-19
c60 77 Vss 9.32916e-19
c61 72 Vss 0.00720976f
c62 67 Vss 0.00368523f
c63 62 Vss 0.0024107f
c64 57 Vss 0.00389164f
c65 54 Vss 7.92361e-19
c66 48 Vss 0.126059f
c67 43 Vss 0.0296049f
c68 39 Vss 2.69463e-19
c69 28 Vss 0.152395f
c70 24 Vss 2.35358e-19
c71 21 Vss 0.169387f
c72 18 Vss 0.0715834f
c73 16 Vss 0.0247918f
c74 10 Vss 0.0674191f
c75 7 Vss 0.219218f
c76 4 Vss 0.08397f
r77 81 85 0.653045
r78 62 77 1.16709
r79 62 85 4.9014
r80 57 72 1.16709
r81 57 81 8.169
r82 51 67 1.16709
r83 51 54 0.0364688
r84 47 72 0.262036
r85 47 48 2.334
r86 44 47 2.20433
r87 39 77 0.404964
r88 33 48 0.00605528
r89 31 44 0.00605528
r90 29 43 0.494161
r91 28 30 0.652036
r92 28 29 4.84305
r93 25 43 0.128424
r94 24 67 0.0476429
r95 22 24 0.326018
r96 22 24 0.1167
r97 21 43 0.494161
r98 21 24 6.7686
r99 18 67 0.357321
r100 16 24 0.326018
r101 16 18 0.40845
r102 10 39 2.04225
r103 7 33 2.5674
r104 7 31 2.5674
r105 7 30 2.5674
r106 4 25 2.5674
r107 2 18 2.15895
.ends

.subckt PM_G4_XOR2_N1_NET1 2 7 10 31 35 44 49 58 76 Vss
c41 76 Vss 3.74063e-19
c42 58 Vss 0.00478125f
c43 49 Vss 0.00566108f
c44 44 Vss 0.0016591f
c45 35 Vss 0.102425f
c46 31 Vss 0.123619f
c47 10 Vss 0.181762f
c48 7 Vss 0.270505f
c49 2 Vss 0.00157712f
r50 72 76 0.653045
r51 49 58 1.16709
r52 49 76 12.9148
r53 44 72 2.08393
r54 33 35 1.70187
r55 30 58 0.262036
r56 30 31 2.20433
r57 27 30 2.334
r58 25 35 0.17282
r59 24 31 0.00605528
r60 21 33 0.17282
r61 18 27 0.00605528
r62 10 21 5.77665
r63 7 25 4.4346
r64 7 24 2.5674
r65 7 18 2.5674
r66 2 44 1.16709
.ends

.subckt PM_G4_XOR2_N1_NET2 2 6 9 21 22 32 33 42 47 56 74 Vss
c46 74 Vss 3.38305e-19
c47 56 Vss 0.00607606f
c48 47 Vss 0.00639628f
c49 42 Vss 0.00204719f
c50 33 Vss 0.126868f
c51 22 Vss 0.0327936f
c52 21 Vss 0.172441f
c53 9 Vss 0.361367f
c54 6 Vss 0.09048f
c55 2 Vss 0.00157712f
r56 70 74 0.660011
r57 47 56 1.16709
r58 47 74 11.3611
r59 42 70 1.95889
r60 32 56 0.262036
r61 32 33 2.26917
r62 29 32 2.26917
r63 26 33 0.00605528
r64 24 29 0.00605528
r65 21 23 0.652036
r66 21 22 4.84305
r67 18 22 0.652036
r68 9 26 2.5674
r69 9 24 2.5674
r70 9 23 7.4688
r71 6 18 2.97585
r72 2 42 1.16709
.ends

.subckt PM_G4_XOR2_N1_B 2 4 7 10 19 20 28 31 36 47 49 52 55 58 61 Vss
c39 61 Vss 0.0281877f
c40 58 Vss 0.00108886f
c41 52 Vss 0.0966253f
c42 49 Vss 0.0299431f
c43 47 Vss 0.131329f
c44 36 Vss 0.043285f
c45 31 Vss 2.35358e-19
c46 28 Vss 0.117434f
c47 20 Vss 0.03478f
c48 19 Vss 0.169387f
c49 10 Vss 0.155214f
c50 7 Vss 0.215531f
c51 4 Vss 0.0714224f
c52 2 Vss 0.083716f
r53 58 61 1.16709
r54 55 58 0.0729375
r55 50 52 2.04225
r56 45 47 4.53833
r57 40 47 0.00605528
r58 37 52 0.0685365
r59 36 50 0.0685365
r60 35 49 0.494161
r61 35 36 1.69215
r62 33 49 0.494161
r63 32 45 0.00605528
r64 31 61 0.181909
r65 29 61 0.494161
r66 29 31 0.1167
r67 28 49 0.128424
r68 28 31 4.72635
r69 23 61 0.128424
r70 23 61 0.40845
r71 22 61 0.181909
r72 20 22 6.7686
r73 19 61 0.494161
r74 19 22 0.1167
r75 16 20 0.652036
r76 10 37 5.0181
r77 7 40 2.5674
r78 7 33 2.5674
r79 7 32 2.5674
r80 4 61 2.15895
r81 2 16 2.5674
.ends

.subckt PM_G4_XOR2_N1_Z 2 4 30 33 Vss
c26 30 Vss 0.00301247f
c27 4 Vss 0.00253802f
c28 2 Vss 0.00148239f
r29 33 35 3.12589
r30 30 33 5.16814
r31 4 35 1.16709
r32 2 30 1.16709
.ends

.subckt G4_XOR2_N1  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI1.X0 N_NET1_XI1.X0_D N_VDD_XI1.X0_PGD N_B_XI1.X0_CG N_VDD_XI1.X0_PGD
+ N_VSS_XI1.X0_S TIGFET_HPNW4
XI9.X0 N_NET2_XI9.X0_D N_VSS_XI9.X0_PGD N_A_XI9.X0_CG N_VSS_XI9.X0_PGD
+ N_VDD_XI9.X0_S TIGFET_HPNW4
XI10.X0 N_NET1_XI1.X0_D N_VSS_XI10.X0_PGD N_B_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW4
XI3.X0 N_NET2_XI9.X0_D N_VDD_XI3.X0_PGD N_A_XI3.X0_CG N_VDD_XI3.X0_PGD
+ N_VSS_XI3.X0_S TIGFET_HPNW4
XI5.X0 N_Z_XI5.X0_D N_B_XI5.X0_PGD N_NET2_XI5.X0_CG N_B_XI5.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW4
XI8.X0 N_Z_XI8.X0_D N_A_XI8.X0_PGD N_B_XI8.X0_CG N_A_XI8.X0_PGD N_VSS_XI3.X0_S
+ TIGFET_HPNW4
XI11.X0 N_Z_XI5.X0_D N_NET1_XI11.X0_PGD N_A_XI11.X0_CG N_NET1_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW4
XI7.X0 N_Z_XI8.X0_D N_NET2_XI7.X0_PGD N_NET1_XI7.X0_CG N_NET2_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW4
*
x_PM_G4_XOR2_N1_VSS N_VSS_XI1.X0_S N_VSS_XI9.X0_PGD N_VSS_XI10.X0_PGD
+ N_VSS_XI3.X0_S N_VSS_XI7.X0_S N_VSS_c_8_p N_VSS_c_23_p N_VSS_c_56_p
+ N_VSS_c_40_p N_VSS_c_7_p N_VSS_c_3_p N_VSS_c_13_p N_VSS_c_30_p N_VSS_c_4_p
+ N_VSS_c_6_p N_VSS_c_14_p N_VSS_c_31_p N_VSS_c_10_p N_VSS_c_11_p N_VSS_c_18_p
+ N_VSS_c_19_p N_VSS_c_26_p N_VSS_c_29_p N_VSS_c_27_p N_VSS_c_62_p N_VSS_c_46_p
+ N_VSS_c_83_p N_VSS_c_12_p N_VSS_c_28_p VSS Vss PM_G4_XOR2_N1_VSS
x_PM_G4_XOR2_N1_VDD N_VDD_XI1.X0_PGD N_VDD_XI9.X0_S N_VDD_XI10.X0_S
+ N_VDD_XI3.X0_PGD N_VDD_XI11.X0_S N_VDD_c_112_n N_VDD_c_163_p N_VDD_c_113_n
+ N_VDD_c_114_n N_VDD_c_118_n N_VDD_c_121_n N_VDD_c_124_n N_VDD_c_125_n
+ N_VDD_c_127_n N_VDD_c_134_n N_VDD_c_135_n N_VDD_c_137_n N_VDD_c_141_n
+ N_VDD_c_144_n N_VDD_c_168_p N_VDD_c_149_n N_VDD_c_182_p N_VDD_c_152_n
+ N_VDD_c_153_n VDD N_VDD_c_154_n N_VDD_c_156_n Vss PM_G4_XOR2_N1_VDD
x_PM_G4_XOR2_N1_A N_A_XI9.X0_CG N_A_XI3.X0_CG N_A_XI8.X0_PGD N_A_XI11.X0_CG
+ N_A_c_212_n N_A_c_213_n N_A_c_215_n N_A_c_216_n N_A_c_246_p N_A_c_231_n A
+ N_A_c_219_n N_A_c_223_n N_A_c_224_n N_A_c_239_n N_A_c_242_p N_A_c_240_n Vss
+ PM_G4_XOR2_N1_A
x_PM_G4_XOR2_N1_NET1 N_NET1_XI1.X0_D N_NET1_XI11.X0_PGD N_NET1_XI7.X0_CG
+ N_NET1_c_282_n N_NET1_c_302_p N_NET1_c_273_n N_NET1_c_276_n N_NET1_c_289_n
+ N_NET1_c_277_n Vss PM_G4_XOR2_N1_NET1
x_PM_G4_XOR2_N1_NET2 N_NET2_XI9.X0_D N_NET2_XI5.X0_CG N_NET2_XI7.X0_PGD
+ N_NET2_c_333_n N_NET2_c_352_p N_NET2_c_334_n N_NET2_c_335_n N_NET2_c_314_n
+ N_NET2_c_318_n N_NET2_c_338_n N_NET2_c_321_n Vss PM_G4_XOR2_N1_NET2
x_PM_G4_XOR2_N1_B N_B_XI1.X0_CG N_B_XI10.X0_CG N_B_XI5.X0_PGD N_B_XI8.X0_CG
+ N_B_c_360_n N_B_c_381_n N_B_c_362_n N_B_c_363_n N_B_c_392_n N_B_c_364_n
+ N_B_c_393_n N_B_c_383_n B N_B_c_365_n N_B_c_367_n Vss PM_G4_XOR2_N1_B
x_PM_G4_XOR2_N1_Z N_Z_XI5.X0_D N_Z_XI8.X0_D N_Z_c_401_n Z Vss PM_G4_XOR2_N1_Z
cc_1 N_VSS_XI9.X0_PGD N_VDD_XI1.X0_PGD 2.77144e-19
cc_2 N_VSS_XI10.X0_PGD N_VDD_XI1.X0_PGD 0.00167677f
cc_3 N_VSS_c_3_p N_VDD_XI9.X0_S 2.05974e-19
cc_4 N_VSS_c_4_p N_VDD_XI10.X0_S 2.02468e-19
cc_5 N_VSS_XI9.X0_PGD N_VDD_XI3.X0_PGD 0.00169392f
cc_6 N_VSS_c_6_p N_VDD_XI11.X0_S 2.02468e-19
cc_7 N_VSS_c_7_p N_VDD_c_112_n 0.00167677f
cc_8 N_VSS_c_8_p N_VDD_c_113_n 0.00169392f
cc_9 N_VSS_c_3_p N_VDD_c_114_n 0.00187494f
cc_10 N_VSS_c_10_p N_VDD_c_114_n 0.00305883f
cc_11 N_VSS_c_11_p N_VDD_c_114_n 0.00593001f
cc_12 N_VSS_c_12_p N_VDD_c_114_n 8.91588e-19
cc_13 N_VSS_c_13_p N_VDD_c_118_n 4.43871e-19
cc_14 N_VSS_c_14_p N_VDD_c_118_n 3.66936e-19
cc_15 N_VSS_c_11_p N_VDD_c_118_n 0.0030181f
cc_16 N_VSS_XI1.X0_S N_VDD_c_121_n 3.7884e-19
cc_17 N_VSS_c_3_p N_VDD_c_121_n 4.73473e-19
cc_18 N_VSS_c_18_p N_VDD_c_121_n 0.00352628f
cc_19 N_VSS_c_19_p N_VDD_c_124_n 0.0010586f
cc_20 N_VSS_XI1.X0_S N_VDD_c_125_n 2.02468e-19
cc_21 N_VSS_c_3_p N_VDD_c_125_n 8.57018e-19
cc_22 N_VSS_c_8_p N_VDD_c_127_n 3.60588e-19
cc_23 N_VSS_c_23_p N_VDD_c_127_n 3.60588e-19
cc_24 N_VSS_c_13_p N_VDD_c_127_n 0.00141228f
cc_25 N_VSS_c_14_p N_VDD_c_127_n 0.00112249f
cc_26 N_VSS_c_26_p N_VDD_c_127_n 0.00343125f
cc_27 N_VSS_c_27_p N_VDD_c_127_n 0.0059942f
cc_28 N_VSS_c_28_p N_VDD_c_127_n 7.74609e-19
cc_29 N_VSS_c_29_p N_VDD_c_134_n 0.00107456f
cc_30 N_VSS_c_30_p N_VDD_c_135_n 9.22488e-19
cc_31 N_VSS_c_31_p N_VDD_c_135_n 3.82294e-19
cc_32 N_VSS_c_7_p N_VDD_c_137_n 3.60588e-19
cc_33 N_VSS_c_30_p N_VDD_c_137_n 0.00161703f
cc_34 N_VSS_c_31_p N_VDD_c_137_n 2.03837e-19
cc_35 N_VSS_c_18_p N_VDD_c_137_n 0.00605426f
cc_36 N_VSS_c_13_p N_VDD_c_141_n 9.25616e-19
cc_37 N_VSS_c_4_p N_VDD_c_141_n 9.18823e-19
cc_38 N_VSS_c_14_p N_VDD_c_141_n 3.99794e-19
cc_39 N_VSS_XI3.X0_S N_VDD_c_144_n 2.21516e-19
cc_40 N_VSS_c_40_p N_VDD_c_144_n 2.69489e-19
cc_41 N_VSS_c_30_p N_VDD_c_144_n 0.0023129f
cc_42 N_VSS_c_4_p N_VDD_c_144_n 2.43341e-19
cc_43 N_VSS_c_31_p N_VDD_c_144_n 9.55109e-19
cc_44 N_VSS_XI7.X0_S N_VDD_c_149_n 2.02468e-19
cc_45 N_VSS_c_6_p N_VDD_c_149_n 2.98086e-19
cc_46 N_VSS_c_46_p N_VDD_c_149_n 0.00130737f
cc_47 N_VSS_c_11_p N_VDD_c_152_n 9.23211e-19
cc_48 N_VSS_c_18_p N_VDD_c_153_n 0.0010761f
cc_49 N_VSS_c_30_p N_VDD_c_154_n 3.48267e-19
cc_50 N_VSS_c_31_p N_VDD_c_154_n 8.0279e-19
cc_51 N_VSS_c_13_p N_VDD_c_156_n 3.48267e-19
cc_52 N_VSS_c_14_p N_VDD_c_156_n 8.07896e-19
cc_53 N_VSS_c_14_p N_A_c_212_n 0.00234108f
cc_54 N_VSS_XI9.X0_PGD N_A_c_213_n 3.99472e-19
cc_55 N_VSS_XI10.X0_PGD N_A_c_213_n 2.20169e-19
cc_56 N_VSS_c_56_p N_A_c_215_n 9.41527e-19
cc_57 N_VSS_XI10.X0_PGD N_A_c_216_n 2.20169e-19
cc_58 N_VSS_c_13_p A 5.59945e-19
cc_59 N_VSS_c_14_p A 4.56568e-19
cc_60 N_VSS_c_4_p N_A_c_219_n 0.00506909f
cc_61 N_VSS_c_11_p N_A_c_219_n 6.18143e-19
cc_62 N_VSS_c_62_p N_A_c_219_n 0.00198136f
cc_63 N_VSS_c_46_p N_A_c_219_n 2.97351e-19
cc_64 N_VSS_c_62_p N_A_c_223_n 0.00118029f
cc_65 N_VSS_c_13_p N_A_c_224_n 4.56568e-19
cc_66 N_VSS_c_14_p N_A_c_224_n 6.1245e-19
cc_67 N_VSS_XI1.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_68 N_VSS_c_3_p N_NET1_XI1.X0_D 3.48267e-19
cc_69 N_VSS_XI1.X0_S N_NET1_c_273_n 3.48267e-19
cc_70 N_VSS_c_3_p N_NET1_c_273_n 0.00108327f
cc_71 N_VSS_c_18_p N_NET1_c_273_n 3.32126e-19
cc_72 N_VSS_c_30_p N_NET1_c_276_n 0.00167316f
cc_73 N_VSS_c_10_p N_NET1_c_277_n 3.27829e-19
cc_74 N_VSS_c_18_p N_NET1_c_277_n 6.3226e-19
cc_75 N_VSS_XI3.X0_S N_NET2_XI9.X0_D 3.43419e-19
cc_76 N_VSS_c_4_p N_NET2_XI9.X0_D 3.48267e-19
cc_77 N_VSS_XI3.X0_S N_NET2_c_314_n 3.48267e-19
cc_78 N_VSS_c_4_p N_NET2_c_314_n 0.00151106f
cc_79 N_VSS_c_11_p N_NET2_c_314_n 5.08641e-19
cc_80 N_VSS_c_27_p N_NET2_c_314_n 3.31434e-19
cc_81 N_VSS_c_4_p N_NET2_c_318_n 0.00228146f
cc_82 N_VSS_c_62_p N_NET2_c_318_n 0.00565735f
cc_83 N_VSS_c_83_p N_NET2_c_318_n 0.00115259f
cc_84 N_VSS_c_13_p N_NET2_c_321_n 5.79036e-19
cc_85 N_VSS_c_27_p N_NET2_c_321_n 0.00176418f
cc_86 N_VSS_c_31_p N_B_XI10.X0_CG 0.00234108f
cc_87 N_VSS_XI10.X0_PGD N_B_XI5.X0_PGD 0.00176522f
cc_88 N_VSS_XI9.X0_PGD N_B_c_360_n 2.20169e-19
cc_89 N_VSS_XI10.X0_PGD N_B_c_360_n 3.99472e-19
cc_90 N_VSS_XI10.X0_PGD N_B_c_362_n 4.05198e-19
cc_91 N_VSS_c_31_p N_B_c_363_n 9.49637e-19
cc_92 N_VSS_c_40_p N_B_c_364_n 0.00154836f
cc_93 N_VSS_c_30_p N_B_c_365_n 5.01474e-19
cc_94 N_VSS_c_31_p N_B_c_365_n 4.56568e-19
cc_95 N_VSS_c_30_p N_B_c_367_n 4.56568e-19
cc_96 N_VSS_c_31_p N_B_c_367_n 6.1245e-19
cc_97 N_VSS_XI3.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_98 N_VSS_XI7.X0_S N_Z_XI8.X0_D 3.43419e-19
cc_99 N_VSS_c_4_p N_Z_XI8.X0_D 3.48267e-19
cc_100 N_VSS_c_6_p N_Z_XI8.X0_D 3.48267e-19
cc_101 N_VSS_XI3.X0_S N_Z_c_401_n 3.48267e-19
cc_102 N_VSS_XI7.X0_S N_Z_c_401_n 3.48267e-19
cc_103 N_VSS_c_4_p N_Z_c_401_n 4.94062e-19
cc_104 N_VSS_c_6_p N_Z_c_401_n 5.68744e-19
cc_105 N_VSS_c_62_p N_Z_c_401_n 3.25705e-19
cc_106 N_VDD_c_156_n N_A_XI3.X0_CG 9.28877e-19
cc_107 N_VDD_XI3.X0_PGD N_A_XI8.X0_PGD 0.00157721f
cc_108 N_VDD_XI1.X0_PGD N_A_c_213_n 2.20169e-19
cc_109 N_VDD_XI3.X0_PGD N_A_c_213_n 4.04053e-19
cc_110 N_VDD_XI3.X0_PGD N_A_c_216_n 4.05198e-19
cc_111 N_VDD_c_163_p N_A_c_231_n 0.00157721f
cc_112 N_VDD_c_114_n A 3.46645e-19
cc_113 N_VDD_c_135_n A 2.52205e-19
cc_114 N_VDD_c_141_n N_A_c_219_n 5.08705e-19
cc_115 N_VDD_c_156_n N_A_c_219_n 3.5189e-19
cc_116 N_VDD_c_168_p N_A_c_223_n 8.44396e-19
cc_117 N_VDD_c_114_n N_A_c_224_n 4.71537e-19
cc_118 N_VDD_c_154_n N_A_c_224_n 4.4222e-19
cc_119 N_VDD_c_156_n N_A_c_239_n 9.06702e-19
cc_120 N_VDD_c_168_p N_A_c_240_n 0.00102412f
cc_121 N_VDD_XI10.X0_S N_NET1_XI1.X0_D 3.43419e-19
cc_122 N_VDD_c_137_n N_NET1_XI1.X0_D 3.7884e-19
cc_123 N_VDD_c_144_n N_NET1_XI1.X0_D 3.48267e-19
cc_124 N_VDD_c_168_p N_NET1_c_282_n 8.23105e-19
cc_125 N_VDD_XI10.X0_S N_NET1_c_273_n 3.48267e-19
cc_126 N_VDD_c_137_n N_NET1_c_273_n 4.58491e-19
cc_127 N_VDD_c_144_n N_NET1_c_273_n 0.00110118f
cc_128 N_VDD_c_144_n N_NET1_c_276_n 0.00124814f
cc_129 N_VDD_c_168_p N_NET1_c_276_n 0.00341061f
cc_130 N_VDD_c_182_p N_NET1_c_276_n 8.21148e-19
cc_131 N_VDD_c_144_n N_NET1_c_289_n 2.78343e-19
cc_132 N_VDD_c_168_p N_NET1_c_289_n 0.00115624f
cc_133 N_VDD_c_182_p N_NET1_c_289_n 3.70842e-19
cc_134 N_VDD_c_135_n N_NET1_c_277_n 2.90608e-19
cc_135 N_VDD_XI9.X0_S N_NET2_XI9.X0_D 3.67949e-19
cc_136 N_VDD_c_125_n N_NET2_XI9.X0_D 3.72199e-19
cc_137 N_VDD_XI9.X0_S N_NET2_c_314_n 3.9802e-19
cc_138 N_VDD_c_125_n N_NET2_c_314_n 5.226e-19
cc_139 N_VDD_c_127_n N_NET2_c_314_n 5.01863e-19
cc_140 N_VDD_c_141_n N_NET2_c_318_n 2.9893e-19
cc_141 N_VDD_c_114_n N_B_XI1.X0_CG 3.37985e-19
cc_142 N_VDD_c_154_n N_B_XI1.X0_CG 9.28877e-19
cc_143 N_VDD_XI1.X0_PGD N_B_c_360_n 4.04053e-19
cc_144 N_VDD_XI3.X0_PGD N_B_c_360_n 2.20169e-19
cc_145 N_VDD_XI3.X0_PGD N_B_c_362_n 2.20169e-19
cc_146 N_VDD_c_144_n N_B_c_364_n 2.75901e-19
cc_147 N_VDD_c_168_p N_B_c_364_n 9.79508e-19
cc_148 N_VDD_c_141_n N_B_c_365_n 2.10322e-19
cc_149 N_VDD_c_156_n N_B_c_367_n 4.24849e-19
cc_150 N_VDD_XI10.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_151 N_VDD_XI11.X0_S N_Z_XI5.X0_D 3.43419e-19
cc_152 N_VDD_c_144_n N_Z_XI5.X0_D 3.48267e-19
cc_153 N_VDD_c_168_p N_Z_XI5.X0_D 3.7884e-19
cc_154 N_VDD_c_149_n N_Z_XI5.X0_D 3.72199e-19
cc_155 N_VDD_XI10.X0_S N_Z_c_401_n 3.48267e-19
cc_156 N_VDD_XI11.X0_S N_Z_c_401_n 3.48267e-19
cc_157 N_VDD_c_144_n N_Z_c_401_n 7.90262e-19
cc_158 N_VDD_c_168_p N_Z_c_401_n 6.5261e-19
cc_159 N_VDD_c_149_n N_Z_c_401_n 8.53368e-19
cc_160 N_A_XI11.X0_CG N_NET1_XI11.X0_PGD 4.5346e-19
cc_161 N_A_c_242_p N_NET1_XI11.X0_PGD 0.0013363f
cc_162 N_A_c_223_n N_NET1_c_276_n 0.00121138f
cc_163 N_A_c_240_n N_NET1_c_276_n 0.00197573f
cc_164 N_A_XI11.X0_CG N_NET1_c_289_n 0.00234108f
cc_165 N_A_c_246_p N_NET1_c_289_n 0.00110158f
cc_166 N_A_c_242_p N_NET1_c_289_n 0.0014909f
cc_167 N_A_c_242_p N_NET2_XI5.X0_CG 2.18475e-19
cc_168 N_A_XI8.X0_PGD N_NET2_XI7.X0_PGD 0.00161543f
cc_169 N_A_c_216_n N_NET2_XI7.X0_PGD 3.14428e-19
cc_170 N_A_c_242_p N_NET2_XI7.X0_PGD 4.01857e-19
cc_171 N_A_XI8.X0_PGD N_NET2_c_333_n 4.60549e-19
cc_172 N_A_c_246_p N_NET2_c_334_n 2.17364e-19
cc_173 N_A_c_231_n N_NET2_c_335_n 0.00161543f
cc_174 N_A_c_219_n N_NET2_c_318_n 0.00221613f
cc_175 N_A_c_223_n N_NET2_c_318_n 7.30894e-19
cc_176 N_A_c_219_n N_NET2_c_338_n 3.44698e-19
cc_177 N_A_c_239_n N_NET2_c_338_n 9.17176e-19
cc_178 N_A_c_242_p N_NET2_c_338_n 3.34137e-19
cc_179 N_A_c_216_n N_B_XI8.X0_CG 0.003858f
cc_180 N_A_c_239_n N_B_XI8.X0_CG 0.00111269f
cc_181 N_A_c_213_n N_B_c_360_n 0.00504555f
cc_182 N_A_c_224_n N_B_c_381_n 3.67702e-19
cc_183 N_A_c_216_n N_B_c_362_n 0.00373351f
cc_184 N_A_c_216_n N_B_c_383_n 0.00215664f
cc_185 N_A_c_240_n N_B_c_365_n 2.66007e-19
cc_186 N_A_c_213_n N_B_c_367_n 4.25664e-19
cc_187 N_A_c_219_n N_Z_c_401_n 0.00323423f
cc_188 N_A_c_223_n N_Z_c_401_n 0.00319047f
cc_189 N_A_c_242_p N_Z_c_401_n 8.50872e-19
cc_190 N_NET1_c_273_n N_NET2_XI9.X0_D 2.02468e-19
cc_191 N_NET1_XI11.X0_PGD N_NET2_XI5.X0_CG 3.25363e-19
cc_192 N_NET1_c_302_p N_NET2_XI7.X0_PGD 0.00868439f
cc_193 N_NET1_XI11.X0_PGD N_NET2_c_333_n 0.00320236f
cc_194 N_NET1_XI1.X0_D N_NET2_c_314_n 2.02468e-19
cc_195 N_NET1_c_273_n N_NET2_c_314_n 3.48409e-19
cc_196 N_NET1_c_276_n N_NET2_c_318_n 0.00270459f
cc_197 N_NET1_XI7.X0_CG N_NET2_c_338_n 0.00266268f
cc_198 N_NET1_XI11.X0_PGD N_B_XI5.X0_PGD 0.00188194f
cc_199 N_NET1_XI7.X0_CG N_B_XI8.X0_CG 2.72153e-19
cc_200 N_NET1_c_282_n N_B_c_364_n 0.00165596f
cc_201 N_NET1_c_302_p N_B_c_383_n 2.72153e-19
cc_202 N_NET2_XI5.X0_CG N_B_XI5.X0_PGD 0.00233046f
cc_203 N_NET2_c_333_n N_B_XI5.X0_PGD 0.00159876f
cc_204 N_NET2_XI7.X0_PGD N_B_c_392_n 4.0517e-19
cc_205 N_NET2_c_352_p N_B_c_393_n 0.00233046f
cc_206 N_NET2_XI7.X0_PGD N_B_c_383_n 0.00313315f
cc_207 N_NET2_c_352_p N_B_c_383_n 0.00171842f
cc_208 N_NET2_XI7.X0_PGD N_Z_c_401_n 0.0012119f
cc_209 N_NET2_c_333_n N_Z_c_401_n 4.14549e-19
cc_210 N_NET2_c_318_n N_Z_c_401_n 2.62894e-19
cc_211 N_B_c_383_n N_Z_c_401_n 8.74847e-19
*
.ends
*
*
.subckt XOR2_HPNW4 A B Y VDD VSS
xgate (VSS VDD A B Y) G4_XOR2_N1
.ends
*
* File: G5_XOR3_N1.pex.netlist
* Created: Sun Apr 10 19:25:53 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XOR3_N1_VDD 2 5 9 12 14 17 34 35 44 45 54 55 77 79 80 81 84 86 90
+ 93 96 98 102 104 108 114 116 118 120 121 122 128 137 142 Vss
c124 142 Vss 0.00486824f
c125 137 Vss 0.00581297f
c126 128 Vss 0.00564406f
c127 122 Vss 0.0021675f
c128 121 Vss 2.39889e-19
c129 120 Vss 4.91069e-19
c130 119 Vss 4.36646e-19
c131 116 Vss 3.56526e-19
c132 114 Vss 0.00137025f
c133 108 Vss 8.30092e-19
c134 104 Vss 0.00588096f
c135 102 Vss 0.0013924f
c136 98 Vss 0.00493548f
c137 96 Vss 0.00124955f
c138 93 Vss 0.00253806f
c139 90 Vss 0.00359127f
c140 86 Vss 0.0066064f
c141 84 Vss 0.0015095f
c142 81 Vss 8.67096e-19
c143 80 Vss 0.0091443f
c144 79 Vss 0.00867106f
c145 77 Vss 0.00186435f
c146 55 Vss 0.0350971f
c147 54 Vss 0.099468f
c148 45 Vss 0.0346156f
c149 44 Vss 0.1003f
c150 35 Vss 0.0346129f
c151 34 Vss 0.0990563f
c152 17 Vss 0.165917f
c153 14 Vss 0.00210084f
c154 12 Vss 0.00231756f
c155 9 Vss 0.16518f
c156 5 Vss 0.165156f
c157 2 Vss 0.00208065f
r158 112 114 4.83471
r159 108 142 1.16709
r160 106 122 0.128424
r161 106 108 2.16729
r162 105 121 0.494161
r163 104 112 0.652036
r164 104 105 7.46046
r165 102 137 1.16709
r166 100 121 0.128424
r167 100 102 2.16729
r168 99 120 0.494161
r169 98 122 0.494161
r170 98 99 10.3363
r171 94 119 0.0828784
r172 94 96 2.00578
r173 93 120 0.128424
r174 92 119 0.551426
r175 92 93 3.91779
r176 90 128 1.16709
r177 88 119 0.551426
r178 88 90 5.835
r179 87 118 0.326018
r180 86 120 0.494161
r181 86 87 10.1279
r182 82 116 0.0828784
r183 82 84 1.82344
r184 80 121 0.494161
r185 80 81 15.8795
r186 79 118 0.326018
r187 78 116 0.551426
r188 78 79 13.0871
r189 77 116 0.551426
r190 76 81 0.652036
r191 76 77 4.16786
r192 57 142 0.0952857
r193 55 57 1.45875
r194 54 58 0.652036
r195 54 57 1.45875
r196 51 55 0.652036
r197 47 137 0.238214
r198 45 47 1.45875
r199 44 48 0.652036
r200 44 47 1.45875
r201 41 45 0.652036
r202 37 128 0.238214
r203 35 37 1.45875
r204 34 38 0.652036
r205 34 37 1.45875
r206 31 35 0.652036
r207 17 58 2.5674
r208 17 51 2.5674
r209 14 114 1.16709
r210 12 96 1.16709
r211 9 48 2.5674
r212 9 41 2.5674
r213 5 38 2.5674
r214 5 31 2.5674
r215 2 84 1.16709
.ends

.subckt PM_G5_XOR3_N1_C 2 4 6 8 17 20 40 43 47 52 57 62 85 87 96 97 Vss
c59 97 Vss 6.9907e-19
c60 87 Vss 0.00433475f
c61 85 Vss 0.00742725f
c62 62 Vss 0.00258068f
c63 57 Vss 0.00592074f
c64 52 Vss 0.00198267f
c65 47 Vss 7.02443e-19
c66 43 Vss 6.02755e-19
c67 40 Vss 6.7024e-19
c68 20 Vss 0.220565f
c69 17 Vss 0.0783954f
c70 15 Vss 0.0247918f
c71 8 Vss 0.00236553f
c72 4 Vss 0.0830741f
r73 88 97 0.0685365
r74 87 89 0.652036
r75 87 88 10.3363
r76 85 97 0.0685365
r77 85 96 24.7154
r78 52 89 2.16729
r79 47 62 1.16709
r80 47 97 2.08393
r81 43 57 1.16709
r82 43 96 0.531835
r83 40 43 0.0833571
r84 23 57 0.238214
r85 21 23 0.326018
r86 21 23 0.1167
r87 20 24 0.652036
r88 20 23 6.7686
r89 17 23 0.262036
r90 15 23 0.326018
r91 15 17 0.05835
r92 8 52 1.16709
r93 6 62 0.8
r94 4 24 2.5674
r95 2 17 2.50905
.ends

.subckt PM_G5_XOR3_N1_VSS 3 6 11 15 18 34 37 44 45 47 54 55 73 78 83 88 93 98
+ 107 112 121 123 124 125 130 131 136 142 153 154 155 156 Vss
c131 156 Vss 3.75522e-19
c132 155 Vss 3.87529e-19
c133 154 Vss 4.4306e-19
c134 142 Vss 0.00208493f
c135 136 Vss 0.00324551f
c136 131 Vss 8.38057e-19
c137 130 Vss 0.00579302f
c138 125 Vss 8.35119e-19
c139 124 Vss 0.00509021f
c140 123 Vss 0.00330591f
c141 121 Vss 0.00273904f
c142 112 Vss 0.00381998f
c143 107 Vss 0.00405934f
c144 98 Vss 0.00484708f
c145 93 Vss 0.00171362f
c146 88 Vss 5.59372e-19
c147 83 Vss 9.83293e-19
c148 78 Vss 0.00292041f
c149 73 Vss 0.00232164f
c150 55 Vss 0.0338093f
c151 54 Vss 0.0988897f
c152 47 Vss 7.82991e-20
c153 45 Vss 0.0347002f
c154 44 Vss 0.0989329f
c155 37 Vss 6.43685e-20
c156 35 Vss 0.0349827f
c157 34 Vss 0.1003f
c158 18 Vss 0.00259162f
c159 15 Vss 0.163916f
c160 11 Vss 0.167978f
c161 6 Vss 0.00155055f
c162 3 Vss 0.167004f
r163 148 153 1.70882
r164 143 156 0.494161
r165 142 148 0.652036
r166 142 143 7.46046
r167 138 156 0.128424
r168 137 155 0.494161
r169 136 144 0.652036
r170 136 137 7.46046
r171 132 155 0.128424
r172 130 156 0.494161
r173 130 131 15.8795
r174 126 154 0.0828784
r175 124 155 0.494161
r176 124 125 13.0037
r177 123 131 0.652036
r178 122 154 0.551426
r179 122 123 10.4196
r180 121 154 0.551426
r181 120 125 0.652036
r182 120 121 6.83529
r183 93 153 2.87582
r184 88 112 1.16709
r185 88 144 2.16729
r186 83 107 1.16709
r187 83 138 2.16729
r188 78 132 4.83471
r189 73 98 1.16709
r190 73 126 4.33978
r191 57 112 0.238214
r192 55 57 1.45875
r193 54 58 0.652036
r194 54 57 1.45875
r195 51 55 0.652036
r196 47 107 0.0952857
r197 45 47 1.45875
r198 44 48 0.652036
r199 44 47 1.45875
r200 41 45 0.652036
r201 37 98 0.238214
r202 35 37 1.45875
r203 34 38 0.652036
r204 34 37 1.45875
r205 31 35 0.652036
r206 18 93 1.16709
r207 15 58 2.5674
r208 15 51 2.5674
r209 11 48 2.5674
r210 11 41 2.5674
r211 6 78 1.16709
r212 3 38 2.5674
r213 3 31 2.5674
.ends

.subckt PM_G5_XOR3_N1_CI 2 6 8 34 39 44 79 80 82 83 84 89 Vss
c62 95 Vss 1.58755e-19
c63 89 Vss 0.00511711f
c64 84 Vss 1.26921e-19
c65 83 Vss 3.02933e-19
c66 82 Vss 0.0013099f
c67 80 Vss 4.32078e-19
c68 79 Vss 0.00369198f
c69 44 Vss 0.00182014f
c70 39 Vss 0.00109627f
c71 34 Vss 0.00267797f
c72 8 Vss 0.00276539f
c73 6 Vss 0.00212882f
c74 2 Vss 0.00154772f
r75 90 95 0.494161
r76 89 91 0.652036
r77 89 90 10.3363
r78 85 95 0.128424
r79 83 95 0.494161
r80 83 84 1.70882
r81 82 84 0.652036
r82 81 82 5.33486
r83 79 81 0.652036
r84 79 80 18.9638
r85 75 80 0.652036
r86 44 91 1.66714
r87 39 85 1.66714
r88 34 75 4.33457
r89 8 44 1.16709
r90 6 39 1.16709
r91 2 34 1.16709
.ends

.subckt PM_G5_XOR3_N1_A 2 4 7 11 21 24 45 49 51 54 55 56 58 62 63 69 74 Vss
c81 74 Vss 0.00494965f
c82 69 Vss 0.00491712f
c83 63 Vss 7.45325e-19
c84 62 Vss 6.24332e-19
c85 56 Vss 0.00115533f
c86 55 Vss 0.00958405f
c87 54 Vss 0.00423116f
c88 51 Vss 0.00507608f
c89 49 Vss 0.135015f
c90 45 Vss 0.125273f
c91 24 Vss 0.213865f
c92 21 Vss 0.0724995f
c93 19 Vss 0.0247918f
c94 7 Vss 1.00758f
c95 4 Vss 0.0850321f
r96 66 74 1.16709
r97 63 66 0.750214
r98 61 69 1.16709
r99 61 62 0.513084
r100 58 61 0.0614211
r101 55 63 0.0685365
r102 55 56 10.4613
r103 53 56 0.652036
r104 53 54 8.66914
r105 51 54 0.652036
r106 51 62 10.2113
r107 47 49 4.53833
r108 44 74 0.262036
r109 44 45 2.26917
r110 41 44 2.26917
r111 36 49 0.00605528
r112 35 45 0.00605528
r113 32 47 0.00605528
r114 31 41 0.00605528
r115 27 69 0.0952857
r116 25 27 0.326018
r117 25 27 0.1167
r118 24 28 0.652036
r119 24 27 6.7686
r120 21 27 0.3335
r121 19 27 0.326018
r122 19 21 0.2334
r123 11 36 2.5674
r124 11 32 2.5674
r125 7 11 12.837
r126 7 35 2.5674
r127 7 11 12.837
r128 7 31 2.5674
r129 4 28 2.5674
r130 2 21 2.334
.ends

.subckt PM_G5_XOR3_N1_BI 2 6 8 18 21 32 37 42 52 57 66 72 73 Vss
c61 73 Vss 1.47395e-19
c62 72 Vss 8.14419e-19
c63 66 Vss 0.00107279f
c64 57 Vss 0.00255458f
c65 52 Vss 0.00234753f
c66 42 Vss 0.00105993f
c67 37 Vss 0.001668f
c68 32 Vss 0.00236426f
c69 21 Vss 0.0573997f
c70 6 Vss 0.0573997f
c71 2 Vss 0.0015046f
r72 72 73 0.655813
r73 71 72 3.501
r74 66 71 0.655813
r75 42 57 1.16709
r76 42 73 2.00578
r77 37 52 1.16709
r78 37 77 12.0712
r79 37 66 2.00578
r80 32 49 1.16709
r81 32 77 2.08393
r82 21 57 0.50025
r83 18 52 0.50025
r84 8 21 1.80885
r85 6 18 1.80885
r86 2 49 0.1
.ends

.subckt PM_G5_XOR3_N1_AI 2 7 11 31 36 37 46 51 60 70 72 82 Vss
c55 82 Vss 2.57983e-19
c56 72 Vss 0.00283715f
c57 70 Vss 0.00386641f
c58 60 Vss 0.00539669f
c59 51 Vss 0.00147157f
c60 46 Vss 0.00243924f
c61 37 Vss 0.127837f
c62 36 Vss 6.45995e-20
c63 31 Vss 0.128147f
c64 7 Vss 0.997493f
c65 2 Vss 0.0015046f
r66 78 82 0.652036
r67 72 82 8.96089
r68 70 74 0.652036
r69 70 72 4.20954
r70 60 63 0.1
r71 51 63 1.16709
r72 51 74 1.83386
r73 46 78 4.58464
r74 36 60 0.262036
r75 36 37 2.334
r76 33 36 2.20433
r77 29 31 4.53833
r78 26 37 0.00605528
r79 25 31 0.00605528
r80 22 33 0.00605528
r81 21 29 0.00605528
r82 11 26 2.5674
r83 11 22 2.5674
r84 7 11 12.837
r85 7 25 2.5674
r86 7 11 12.837
r87 7 21 2.5674
r88 2 46 1.16709
.ends

.subckt PM_G5_XOR3_N1_B 2 4 6 8 16 17 24 26 33 38 42 45 50 55 60 65 73 74 80 86
+ 91 92 Vss
c91 92 Vss 1.10364e-19
c92 91 Vss 9.61135e-19
c93 86 Vss 5.98353e-19
c94 80 Vss 8.23772e-19
c95 74 Vss 5.75465e-19
c96 73 Vss 0.00321909f
c97 65 Vss 0.00250661f
c98 60 Vss 0.00207758f
c99 55 Vss 0.00386058f
c100 50 Vss 0.00113661f
c101 45 Vss 4.31637e-19
c102 42 Vss 4.09773e-19
c103 38 Vss 5.37175e-19
c104 33 Vss 6.95992e-20
c105 26 Vss 0.0573997f
c106 24 Vss 7.82991e-20
c107 20 Vss 0.0247918f
c108 17 Vss 0.0338376f
c109 16 Vss 0.183114f
c110 8 Vss 0.0573997f
c111 4 Vss 0.0714013f
c112 2 Vss 0.0826046f
r113 90 92 0.65228
r114 90 91 3.46076
r115 86 91 0.65228
r116 73 80 0.0685365
r117 73 74 10.3363
r118 69 74 0.652036
r119 50 65 1.16709
r120 50 92 2.1395
r121 45 60 1.16709
r122 45 86 2.1006
r123 45 80 2.08393
r124 38 55 1.16709
r125 38 69 2.16729
r126 38 42 0.0729375
r127 36 55 0.0476429
r128 33 65 0.50025
r129 26 60 0.50025
r130 24 55 0.357321
r131 20 36 0.326018
r132 20 24 0.40845
r133 17 36 6.7686
r134 16 36 0.326018
r135 16 36 0.1167
r136 13 17 0.652036
r137 8 33 1.80885
r138 6 26 1.80885
r139 4 24 2.15895
r140 2 13 2.5674
.ends

.subckt PM_G5_XOR3_N1_Z 2 4 30 33 Vss
c30 30 Vss 0.00324462f
c31 4 Vss 0.00153036f
c32 2 Vss 0.00166246f
r33 33 35 4.50129
r34 30 33 4.668
r35 4 35 1.16709
r36 2 30 1.16709
.ends

.subckt G5_XOR3_N1  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI10.X0 N_CI_XI10.X0_D N_VSS_XI10.X0_PGD N_C_XI10.X0_CG N_VSS_XI10.X0_PGD
+ N_VDD_XI10.X0_S TIGFET_HPNW4
XI9.X0 N_CI_XI10.X0_D N_VDD_XI9.X0_PGD N_C_XI9.X0_CG N_VDD_XI9.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI5.X0 N_BI_XI5.X0_D N_VDD_XI5.X0_PGD N_B_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_VSS_XI9.X0_S TIGFET_HPNW4
XI8.X0 N_AI_XI8.X0_D N_VSS_XI8.X0_PGD N_A_XI8.X0_CG N_VSS_XI8.X0_PGD
+ N_VDD_XI8.X0_S TIGFET_HPNW4
XI6.X0 N_BI_XI5.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW4
XI7.X0 N_AI_XI8.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGD
+ N_VSS_XI7.X0_S TIGFET_HPNW4
XI2.X0 N_Z_XI2.X0_D N_AI_XI2.X0_PGD N_BI_XI2.X0_CG N_AI_XI2.X0_PGD N_C_XI2.X0_S
+ TIGFET_HPNW4
XI4.X0 N_Z_XI4.X0_D N_AI_XI4.X0_PGD N_B_XI4.X0_CG N_AI_XI4.X0_PGD N_CI_XI4.X0_S
+ TIGFET_HPNW4
XI3.X0 N_Z_XI2.X0_D N_A_XI3.X0_PGD N_B_XI3.X0_CG N_A_XI3.X0_PGD N_C_XI3.X0_S
+ TIGFET_HPNW4
XI1.X0 N_Z_XI4.X0_D N_A_XI1.X0_PGD N_BI_XI1.X0_CG N_A_XI1.X0_PGD N_CI_XI1.X0_S
+ TIGFET_HPNW4
*
x_PM_G5_XOR3_N1_VDD N_VDD_XI10.X0_S N_VDD_XI9.X0_PGD N_VDD_XI5.X0_PGD
+ N_VDD_XI8.X0_S N_VDD_XI6.X0_S N_VDD_XI7.X0_PGD N_VDD_c_121_p N_VDD_c_20_p
+ N_VDD_c_25_p N_VDD_c_4_p N_VDD_c_109_p N_VDD_c_21_p N_VDD_c_6_p N_VDD_c_27_p
+ N_VDD_c_5_p N_VDD_c_64_p N_VDD_c_29_p N_VDD_c_30_p N_VDD_c_31_p N_VDD_c_37_p
+ N_VDD_c_34_p N_VDD_c_22_p N_VDD_c_11_p N_VDD_c_26_p N_VDD_c_39_p N_VDD_c_12_p
+ N_VDD_c_60_p VDD N_VDD_c_68_p N_VDD_c_72_p N_VDD_c_19_p N_VDD_c_2_p
+ N_VDD_c_44_p N_VDD_c_40_p Vss PM_G5_XOR3_N1_VDD
x_PM_G5_XOR3_N1_C N_C_XI10.X0_CG N_C_XI9.X0_CG N_C_XI2.X0_S N_C_XI3.X0_S
+ N_C_c_144_p N_C_c_127_n C N_C_c_140_p N_C_c_157_p N_C_c_179_p N_C_c_132_n
+ N_C_c_134_n N_C_c_135_n N_C_c_156_p N_C_c_141_p N_C_c_160_p Vss
+ PM_G5_XOR3_N1_C
x_PM_G5_XOR3_N1_VSS N_VSS_XI10.X0_PGD N_VSS_XI9.X0_S N_VSS_XI8.X0_PGD
+ N_VSS_XI6.X0_PGD N_VSS_XI7.X0_S N_VSS_c_191_n N_VSS_c_250_n N_VSS_c_192_n
+ N_VSS_c_194_n N_VSS_c_288_p N_VSS_c_195_n N_VSS_c_196_n N_VSS_c_198_n
+ N_VSS_c_204_n N_VSS_c_208_n N_VSS_c_212_n N_VSS_c_216_n N_VSS_c_218_n
+ N_VSS_c_221_n N_VSS_c_225_n N_VSS_c_229_n N_VSS_c_232_n N_VSS_c_234_n
+ N_VSS_c_235_n N_VSS_c_236_n N_VSS_c_240_n N_VSS_c_241_n N_VSS_c_244_n VSS
+ N_VSS_c_246_n N_VSS_c_247_n N_VSS_c_248_n Vss PM_G5_XOR3_N1_VSS
x_PM_G5_XOR3_N1_CI N_CI_XI10.X0_D N_CI_XI4.X0_S N_CI_XI1.X0_S N_CI_c_317_n
+ N_CI_c_333_n N_CI_c_373_p N_CI_c_321_n N_CI_c_337_n N_CI_c_339_n N_CI_c_347_p
+ N_CI_c_356_p N_CI_c_325_n Vss PM_G5_XOR3_N1_CI
x_PM_G5_XOR3_N1_A N_A_XI8.X0_CG N_A_XI7.X0_CG N_A_XI3.X0_PGD N_A_XI1.X0_PGD
+ N_A_c_402_n N_A_c_378_n N_A_c_428_p N_A_c_430_p N_A_c_379_n N_A_c_387_n
+ N_A_c_396_n N_A_c_388_n A N_A_c_389_n N_A_c_401_n N_A_c_390_n N_A_c_434_p Vss
+ PM_G5_XOR3_N1_A
x_PM_G5_XOR3_N1_BI N_BI_XI5.X0_D N_BI_XI2.X0_CG N_BI_XI1.X0_CG N_BI_c_480_n
+ N_BI_c_481_n N_BI_c_460_n N_BI_c_464_n N_BI_c_478_n N_BI_c_486_n N_BI_c_487_n
+ N_BI_c_467_n N_BI_c_506_p N_BI_c_479_n Vss PM_G5_XOR3_N1_BI
x_PM_G5_XOR3_N1_AI N_AI_XI8.X0_D N_AI_XI2.X0_PGD N_AI_XI4.X0_PGD N_AI_c_532_n
+ N_AI_c_566_p N_AI_c_522_n N_AI_c_523_n N_AI_c_537_n N_AI_c_527_n N_AI_c_528_n
+ N_AI_c_529_n N_AI_c_540_n Vss PM_G5_XOR3_N1_AI
x_PM_G5_XOR3_N1_B N_B_XI5.X0_CG N_B_XI6.X0_CG N_B_XI4.X0_CG N_B_XI3.X0_CG
+ N_B_c_576_n N_B_c_578_n N_B_c_590_n N_B_c_648_n N_B_c_611_n N_B_c_579_n B
+ N_B_c_615_n N_B_c_583_n N_B_c_580_n N_B_c_620_n N_B_c_621_n N_B_c_581_n
+ N_B_c_602_n N_B_c_603_n N_B_c_585_n N_B_c_645_n N_B_c_586_n Vss
+ PM_G5_XOR3_N1_B
x_PM_G5_XOR3_N1_Z N_Z_XI2.X0_D N_Z_XI4.X0_D N_Z_c_669_n Z Vss PM_G5_XOR3_N1_Z
cc_1 N_VDD_XI5.X0_PGD N_C_XI9.X0_CG 9.6041e-19
cc_2 N_VDD_c_2_p N_C_XI9.X0_CG 8.03148e-19
cc_3 N_VDD_XI9.X0_PGD N_C_c_127_n 4.16623e-19
cc_4 N_VDD_c_4_p N_C_c_127_n 9.6041e-19
cc_5 N_VDD_c_5_p N_C_c_127_n 0.00125128f
cc_6 N_VDD_c_6_p C 4.36744e-19
cc_7 N_VDD_c_5_p C 0.00161703f
cc_8 N_VDD_c_6_p N_C_c_132_n 3.66936e-19
cc_9 N_VDD_c_5_p N_C_c_132_n 2.84956e-19
cc_10 N_VDD_XI6.X0_S N_C_c_134_n 3.43419e-19
cc_11 N_VDD_c_11_p N_C_c_135_n 4.67477e-19
cc_12 N_VDD_c_12_p N_C_c_135_n 7.7658e-19
cc_13 N_VDD_XI9.X0_PGD N_VSS_XI10.X0_PGD 0.00173038f
cc_14 N_VDD_c_5_p N_VSS_XI9.X0_S 3.7884e-19
cc_15 N_VDD_XI5.X0_PGD N_VSS_XI8.X0_PGD 2.27468e-19
cc_16 N_VDD_XI7.X0_PGD N_VSS_XI8.X0_PGD 0.00172148f
cc_17 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.0017188f
cc_18 N_VDD_XI7.X0_PGD N_VSS_XI6.X0_PGD 2.1536e-19
cc_19 N_VDD_c_19_p N_VSS_XI7.X0_S 4.04413e-19
cc_20 N_VDD_c_20_p N_VSS_c_191_n 0.00173038f
cc_21 N_VDD_c_21_p N_VSS_c_192_n 0.00172148f
cc_22 N_VDD_c_22_p N_VSS_c_192_n 2.51785e-19
cc_23 N_VDD_c_22_p N_VSS_c_194_n 3.71017e-19
cc_24 N_VDD_c_12_p N_VSS_c_195_n 2.35445e-19
cc_25 N_VDD_c_25_p N_VSS_c_196_n 0.0017188f
cc_26 N_VDD_c_26_p N_VSS_c_196_n 2.74208e-19
cc_27 N_VDD_c_27_p N_VSS_c_198_n 4.32468e-19
cc_28 N_VDD_c_5_p N_VSS_c_198_n 4.60511e-19
cc_29 N_VDD_c_29_p N_VSS_c_198_n 0.00130521f
cc_30 N_VDD_c_30_p N_VSS_c_198_n 4.5978e-19
cc_31 N_VDD_c_31_p N_VSS_c_198_n 3.98949e-19
cc_32 N_VDD_c_2_p N_VSS_c_198_n 3.48267e-19
cc_33 N_VDD_c_5_p N_VSS_c_204_n 4.58491e-19
cc_34 N_VDD_c_34_p N_VSS_c_204_n 2.25587e-19
cc_35 N_VDD_c_11_p N_VSS_c_204_n 7.77634e-19
cc_36 N_VDD_c_12_p N_VSS_c_204_n 3.28649e-19
cc_37 N_VDD_c_37_p N_VSS_c_208_n 4.0876e-19
cc_38 N_VDD_c_22_p N_VSS_c_208_n 0.00141228f
cc_39 N_VDD_c_39_p N_VSS_c_208_n 8.73606e-19
cc_40 N_VDD_c_40_p N_VSS_c_208_n 3.48267e-19
cc_41 N_VDD_c_11_p N_VSS_c_212_n 6.87451e-19
cc_42 N_VDD_c_26_p N_VSS_c_212_n 0.00141228f
cc_43 N_VDD_c_12_p N_VSS_c_212_n 0.00254823f
cc_44 N_VDD_c_44_p N_VSS_c_212_n 3.48267e-19
cc_45 N_VDD_c_39_p N_VSS_c_216_n 7.30795e-19
cc_46 N_VDD_c_19_p N_VSS_c_216_n 5.00098e-19
cc_47 N_VDD_c_27_p N_VSS_c_218_n 4.41003e-19
cc_48 N_VDD_c_31_p N_VSS_c_218_n 3.89161e-19
cc_49 N_VDD_c_2_p N_VSS_c_218_n 7.99831e-19
cc_50 N_VDD_c_37_p N_VSS_c_221_n 3.48267e-19
cc_51 N_VDD_c_22_p N_VSS_c_221_n 0.00112249f
cc_52 N_VDD_c_39_p N_VSS_c_221_n 3.99794e-19
cc_53 N_VDD_c_40_p N_VSS_c_221_n 8.07559e-19
cc_54 N_VDD_c_11_p N_VSS_c_225_n 3.82294e-19
cc_55 N_VDD_c_26_p N_VSS_c_225_n 0.00112249f
cc_56 N_VDD_c_12_p N_VSS_c_225_n 9.55109e-19
cc_57 N_VDD_c_44_p N_VSS_c_225_n 8.01441e-19
cc_58 N_VDD_c_6_p N_VSS_c_229_n 0.003116f
cc_59 N_VDD_c_27_p N_VSS_c_229_n 7.60301e-19
cc_60 N_VDD_c_60_p N_VSS_c_229_n 0.0010705f
cc_61 N_VDD_c_27_p N_VSS_c_232_n 0.00754268f
cc_62 N_VDD_c_31_p N_VSS_c_232_n 9.72927e-19
cc_63 N_VDD_c_5_p N_VSS_c_234_n 0.00967241f
cc_64 N_VDD_c_64_p N_VSS_c_235_n 0.00107121f
cc_65 N_VDD_c_30_p N_VSS_c_236_n 0.0081111f
cc_66 N_VDD_c_34_p N_VSS_c_236_n 7.52646e-19
cc_67 N_VDD_c_22_p N_VSS_c_236_n 0.00375883f
cc_68 N_VDD_c_68_p N_VSS_c_236_n 0.0014027f
cc_69 N_VDD_c_27_p N_VSS_c_240_n 0.00107333f
cc_70 N_VDD_c_5_p N_VSS_c_241_n 0.00142828f
cc_71 N_VDD_c_26_p N_VSS_c_241_n 0.00543165f
cc_72 N_VDD_c_72_p N_VSS_c_241_n 0.00106247f
cc_73 N_VDD_c_22_p N_VSS_c_244_n 0.00372698f
cc_74 N_VDD_c_19_p N_VSS_c_244_n 0.00347642f
cc_75 N_VDD_c_27_p N_VSS_c_246_n 0.00112682f
cc_76 N_VDD_c_5_p N_VSS_c_247_n 0.00104966f
cc_77 N_VDD_c_22_p N_VSS_c_248_n 7.74609e-19
cc_78 N_VDD_XI10.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_79 N_VDD_c_29_p N_CI_XI10.X0_D 3.72199e-19
cc_80 N_VDD_XI10.X0_S N_CI_c_317_n 3.48267e-19
cc_81 N_VDD_c_5_p N_CI_c_317_n 5.01863e-19
cc_82 N_VDD_c_29_p N_CI_c_317_n 5.226e-19
cc_83 N_VDD_c_31_p N_CI_c_317_n 4.13481e-19
cc_84 N_VDD_c_31_p N_CI_c_321_n 7.11597e-19
cc_85 N_VDD_c_34_p N_CI_c_321_n 7.78475e-19
cc_86 N_VDD_c_40_p N_A_XI7.X0_CG 0.00119068f
cc_87 N_VDD_XI7.X0_PGD N_A_c_378_n 3.90714e-19
cc_88 N_VDD_XI6.X0_S N_A_c_379_n 2.96819e-19
cc_89 N_VDD_XI7.X0_PGD N_A_c_379_n 2.39692e-19
cc_90 N_VDD_c_22_p N_A_c_379_n 5.16693e-19
cc_91 N_VDD_c_26_p N_A_c_379_n 4.57585e-19
cc_92 N_VDD_c_39_p N_A_c_379_n 5.97577e-19
cc_93 N_VDD_c_12_p N_A_c_379_n 4.47961e-19
cc_94 N_VDD_c_19_p N_A_c_379_n 4.69788e-19
cc_95 N_VDD_c_40_p N_A_c_379_n 4.46731e-19
cc_96 N_VDD_XI6.X0_S N_A_c_387_n 9.18655e-19
cc_97 N_VDD_c_12_p N_A_c_388_n 0.00610545f
cc_98 N_VDD_c_31_p N_A_c_389_n 8.33062e-19
cc_99 N_VDD_c_31_p N_A_c_390_n 6.30148e-19
cc_100 N_VDD_c_44_p N_A_c_390_n 5.39283e-19
cc_101 N_VDD_XI6.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_102 N_VDD_c_12_p N_BI_XI5.X0_D 3.48267e-19
cc_103 N_VDD_XI6.X0_S N_BI_c_460_n 3.48267e-19
cc_104 N_VDD_c_26_p N_BI_c_460_n 4.87462e-19
cc_105 N_VDD_c_12_p N_BI_c_460_n 5.0516e-19
cc_106 N_VDD_XI8.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_107 N_VDD_c_22_p N_AI_XI8.X0_D 4.04413e-19
cc_108 N_VDD_XI7.X0_PGD N_AI_XI2.X0_PGD 2.98495e-19
cc_109 N_VDD_c_109_p N_AI_c_522_n 2.98495e-19
cc_110 N_VDD_XI8.X0_S N_AI_c_523_n 3.48267e-19
cc_111 N_VDD_c_34_p N_AI_c_523_n 4.96286e-19
cc_112 N_VDD_c_22_p N_AI_c_523_n 4.84258e-19
cc_113 N_VDD_c_39_p N_AI_c_523_n 5.74209e-19
cc_114 N_VDD_c_39_p N_AI_c_527_n 2.15672e-19
cc_115 N_VDD_c_19_p N_AI_c_528_n 3.25291e-19
cc_116 N_VDD_c_22_p N_AI_c_529_n 2.81017e-19
cc_117 N_VDD_XI9.X0_PGD N_B_XI5.X0_CG 9.57243e-19
cc_118 N_VDD_c_44_p N_B_XI5.X0_CG 9.74645e-19
cc_119 N_VDD_XI5.X0_PGD N_B_c_576_n 3.9688e-19
cc_120 N_VDD_XI7.X0_PGD N_B_c_576_n 2.07132e-19
cc_121 N_VDD_c_121_p N_B_c_578_n 9.57243e-19
cc_122 N_VDD_c_31_p N_B_c_579_n 6.08224e-19
cc_123 N_VDD_c_40_p N_B_c_580_n 3.47237e-19
cc_124 N_VDD_c_12_p N_B_c_581_n 2.72308e-19
cc_125 N_C_c_127_n N_VSS_XI10.X0_PGD 4.16623e-19
cc_126 N_C_c_132_n N_VSS_c_250_n 6.87259e-19
cc_127 C N_VSS_c_198_n 4.80408e-19
cc_128 N_C_c_140_p N_VSS_c_198_n 3.9981e-19
cc_129 N_C_c_141_p N_VSS_c_198_n 2.54015e-19
cc_130 N_C_c_135_n N_VSS_c_204_n 0.00185659f
cc_131 N_C_c_135_n N_VSS_c_212_n 0.00161389f
cc_132 N_C_c_144_p N_VSS_c_218_n 0.0041277f
cc_133 C N_VSS_c_218_n 4.20453e-19
cc_134 N_C_c_132_n N_VSS_c_218_n 0.00184261f
cc_135 N_C_c_140_p N_VSS_c_229_n 4.01014e-19
cc_136 N_C_c_141_p N_VSS_c_229_n 2.65147e-19
cc_137 C N_VSS_c_234_n 3.52403e-19
cc_138 N_C_c_140_p N_VSS_c_234_n 0.00136475f
cc_139 N_C_c_135_n N_VSS_c_234_n 0.00239048f
cc_140 N_C_c_141_p N_VSS_c_234_n 5.40072e-19
cc_141 N_C_c_135_n N_VSS_c_241_n 0.00182168f
cc_142 N_C_c_135_n N_CI_c_317_n 0.00135409f
cc_143 N_C_c_135_n N_CI_c_321_n 0.0042263f
cc_144 N_C_c_156_p N_CI_c_325_n 6.92841e-19
cc_145 N_C_c_157_p N_A_c_387_n 0.00149093f
cc_146 N_C_c_134_n N_A_c_387_n 8.20481e-19
cc_147 N_C_c_135_n N_A_c_387_n 2.83242e-19
cc_148 N_C_c_160_p N_A_c_387_n 2.26175e-19
cc_149 N_C_c_157_p N_A_c_396_n 0.00194268f
cc_150 N_C_c_134_n N_A_c_396_n 9.18655e-19
cc_151 N_C_c_135_n N_A_c_396_n 4.77334e-19
cc_152 N_C_c_156_p N_A_c_396_n 0.00211066f
cc_153 N_C_c_160_p N_A_c_396_n 6.30333e-19
cc_154 N_C_c_156_p N_A_c_401_n 5.46695e-19
cc_155 N_C_c_135_n N_BI_c_460_n 0.00227671f
cc_156 N_C_c_135_n N_BI_c_464_n 0.00490342f
cc_157 N_C_c_156_p N_BI_c_464_n 0.0015987f
cc_158 N_C_c_160_p N_BI_c_464_n 0.0013513f
cc_159 N_C_c_156_p N_BI_c_467_n 9.86034e-19
cc_160 N_C_c_135_n N_B_c_579_n 2.53746e-19
cc_161 N_C_c_156_p N_B_c_583_n 2.11999e-19
cc_162 N_C_c_157_p N_B_c_581_n 4.78342e-19
cc_163 N_C_c_156_p N_B_c_585_n 5.08651e-19
cc_164 N_C_c_156_p N_B_c_586_n 0.00239488f
cc_165 N_C_XI3.X0_S N_Z_XI2.X0_D 3.43419e-19
cc_166 N_C_c_157_p N_Z_XI2.X0_D 3.48267e-19
cc_167 N_C_c_179_p N_Z_XI2.X0_D 3.48267e-19
cc_168 N_C_c_134_n N_Z_XI2.X0_D 3.43419e-19
cc_169 N_C_XI3.X0_S N_Z_c_669_n 3.48267e-19
cc_170 N_C_c_157_p N_Z_c_669_n 3.23828e-19
cc_171 N_C_c_179_p N_Z_c_669_n 5.71075e-19
cc_172 N_VSS_XI9.X0_S N_CI_XI10.X0_D 3.43419e-19
cc_173 N_VSS_c_204_n N_CI_XI10.X0_D 3.48267e-19
cc_174 N_VSS_XI7.X0_S N_CI_XI4.X0_S 3.43419e-19
cc_175 N_VSS_c_216_n N_CI_XI4.X0_S 3.48267e-19
cc_176 N_VSS_c_198_n N_CI_c_317_n 5.88914e-19
cc_177 N_VSS_c_204_n N_CI_c_317_n 8.48865e-19
cc_178 N_VSS_c_234_n N_CI_c_317_n 3.32126e-19
cc_179 N_VSS_XI7.X0_S N_CI_c_333_n 3.48267e-19
cc_180 N_VSS_c_216_n N_CI_c_333_n 7.99744e-19
cc_181 N_VSS_c_208_n N_CI_c_321_n 3.41088e-19
cc_182 N_VSS_c_244_n N_CI_c_321_n 4.44969e-19
cc_183 N_VSS_c_232_n N_CI_c_337_n 2.78598e-19
cc_184 N_VSS_c_236_n N_CI_c_337_n 0.00159458f
cc_185 N_VSS_c_216_n N_CI_c_339_n 0.00104291f
cc_186 N_VSS_c_221_n N_A_c_402_n 0.00297797f
cc_187 N_VSS_XI8.X0_PGD N_A_c_378_n 3.85826e-19
cc_188 N_VSS_XI7.X0_S N_A_c_379_n 9.18655e-19
cc_189 N_VSS_c_216_n N_A_c_379_n 0.00131738f
cc_190 N_VSS_c_241_n N_A_c_379_n 3.01443e-19
cc_191 N_VSS_c_244_n N_A_c_379_n 5.02211e-19
cc_192 N_VSS_c_208_n N_A_c_389_n 5.62647e-19
cc_193 N_VSS_c_221_n N_A_c_389_n 4.60973e-19
cc_194 N_VSS_c_288_p N_A_c_390_n 9.36847e-19
cc_195 N_VSS_c_208_n N_A_c_390_n 4.56568e-19
cc_196 N_VSS_c_221_n N_A_c_390_n 8.15819e-19
cc_197 N_VSS_XI9.X0_S N_BI_XI5.X0_D 3.43419e-19
cc_198 N_VSS_XI9.X0_S N_BI_c_460_n 3.48267e-19
cc_199 N_VSS_c_204_n N_BI_c_460_n 7.98486e-19
cc_200 N_VSS_c_241_n N_BI_c_460_n 3.20743e-19
cc_201 N_VSS_XI7.X0_S N_AI_XI8.X0_D 3.43419e-19
cc_202 N_VSS_XI6.X0_PGD N_AI_XI2.X0_PGD 2.8463e-19
cc_203 N_VSS_c_195_n N_AI_c_532_n 2.8463e-19
cc_204 N_VSS_XI7.X0_S N_AI_c_523_n 3.48267e-19
cc_205 N_VSS_c_208_n N_AI_c_523_n 0.00108072f
cc_206 N_VSS_c_216_n N_AI_c_523_n 0.00193557f
cc_207 N_VSS_c_244_n N_AI_c_523_n 3.6914e-19
cc_208 N_VSS_c_216_n N_AI_c_537_n 8.20606e-19
cc_209 N_VSS_c_244_n N_AI_c_528_n 9.54335e-19
cc_210 N_VSS_c_244_n N_AI_c_529_n 0.00515467f
cc_211 N_VSS_c_244_n N_AI_c_540_n 0.00185629f
cc_212 N_VSS_c_225_n N_B_XI6.X0_CG 0.00272012f
cc_213 N_VSS_XI8.X0_PGD N_B_c_576_n 2.07132e-19
cc_214 N_VSS_XI6.X0_PGD N_B_c_576_n 3.923e-19
cc_215 N_VSS_c_225_n N_B_c_590_n 0.00130195f
cc_216 N_VSS_c_212_n N_B_c_579_n 7.62066e-19
cc_217 N_VSS_c_212_n B 5.66975e-19
cc_218 N_VSS_c_225_n B 4.56568e-19
cc_219 N_VSS_c_225_n N_B_c_580_n 6.1245e-19
cc_220 N_VSS_c_216_n N_B_c_581_n 6.79536e-19
cc_221 N_CI_c_339_n N_A_c_379_n 6.20926e-19
cc_222 N_CI_c_321_n N_A_c_389_n 0.00116415f
cc_223 N_CI_c_339_n N_A_c_389_n 2.08707e-19
cc_224 N_CI_c_317_n N_BI_c_460_n 5.94242e-19
cc_225 N_CI_c_321_n N_BI_c_460_n 0.00302092f
cc_226 N_CI_c_333_n N_BI_c_464_n 3.50977e-19
cc_227 N_CI_c_321_n N_BI_c_464_n 0.00752744f
cc_228 N_CI_c_347_p N_BI_c_464_n 4.80593e-19
cc_229 N_CI_c_325_n N_BI_c_464_n 5.67893e-19
cc_230 N_CI_c_325_n N_BI_c_478_n 0.00102574f
cc_231 N_CI_c_325_n N_BI_c_479_n 2.55507e-19
cc_232 N_CI_c_321_n N_AI_c_523_n 8.44506e-19
cc_233 N_CI_c_339_n N_AI_c_523_n 0.00100365f
cc_234 N_CI_c_325_n N_AI_c_537_n 0.00169084f
cc_235 N_CI_c_333_n N_AI_c_528_n 8.33462e-19
cc_236 N_CI_c_347_p N_AI_c_528_n 7.14401e-19
cc_237 N_CI_c_356_p N_AI_c_528_n 2.16882e-19
cc_238 N_CI_c_325_n N_AI_c_528_n 5.16616e-19
cc_239 N_CI_c_321_n N_AI_c_529_n 0.00115159f
cc_240 N_CI_c_356_p N_AI_c_529_n 0.00241787f
cc_241 N_CI_c_317_n N_B_c_579_n 2.7112e-19
cc_242 N_CI_c_325_n N_B_c_583_n 7.18914e-19
cc_243 N_CI_c_333_n N_B_c_581_n 8.80932e-19
cc_244 N_CI_c_321_n N_B_c_581_n 0.00348609f
cc_245 N_CI_c_347_p N_B_c_581_n 2.27019e-19
cc_246 N_CI_c_325_n N_B_c_581_n 2.27123e-19
cc_247 N_CI_c_321_n N_B_c_602_n 0.00142048f
cc_248 N_CI_c_339_n N_B_c_603_n 3.62522e-19
cc_249 N_CI_c_339_n N_B_c_585_n 4.56062e-19
cc_250 N_CI_c_325_n N_B_c_585_n 0.00270237f
cc_251 N_CI_XI4.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_252 N_CI_XI1.X0_S N_Z_XI4.X0_D 3.43419e-19
cc_253 N_CI_c_333_n N_Z_XI4.X0_D 3.48267e-19
cc_254 N_CI_c_373_p N_Z_XI4.X0_D 3.48267e-19
cc_255 N_CI_XI4.X0_S N_Z_c_669_n 3.48267e-19
cc_256 N_CI_c_333_n N_Z_c_669_n 5.68744e-19
cc_257 N_CI_c_373_p N_Z_c_669_n 6.06579e-19
cc_258 N_A_c_396_n N_BI_c_480_n 3.17089e-19
cc_259 N_A_XI3.X0_PGD N_BI_c_481_n 8.79767e-19
cc_260 N_A_c_379_n N_BI_c_460_n 4.32688e-19
cc_261 N_A_c_387_n N_BI_c_464_n 9.32646e-19
cc_262 N_A_c_396_n N_BI_c_464_n 5.00869e-19
cc_263 N_A_c_396_n N_BI_c_478_n 3.33012e-19
cc_264 N_A_c_387_n N_BI_c_486_n 3.37713e-19
cc_265 N_A_XI3.X0_PGD N_BI_c_487_n 0.00133285f
cc_266 N_A_c_396_n N_BI_c_467_n 0.00106538f
cc_267 N_A_c_379_n N_AI_XI8.X0_D 9.18655e-19
cc_268 N_A_XI3.X0_PGD N_AI_XI2.X0_PGD 0.0174819f
cc_269 N_A_c_387_n N_AI_XI2.X0_PGD 8.52417e-19
cc_270 N_A_c_428_p N_AI_c_532_n 0.00199595f
cc_271 N_A_c_396_n N_AI_c_532_n 0.00123184f
cc_272 N_A_c_430_p N_AI_c_522_n 0.00202022f
cc_273 N_A_c_379_n N_AI_c_523_n 0.00136181f
cc_274 N_A_c_379_n N_AI_c_529_n 2.67536e-19
cc_275 N_A_XI3.X0_PGD N_B_XI3.X0_CG 8.79767e-19
cc_276 N_A_c_434_p N_B_XI3.X0_CG 0.00237738f
cc_277 N_A_c_378_n N_B_c_576_n 0.0036024f
cc_278 N_A_c_379_n N_B_c_576_n 5.40888e-19
cc_279 N_A_c_390_n N_B_c_578_n 4.08399e-19
cc_280 N_A_c_434_p N_B_c_611_n 0.00115102f
cc_281 N_A_c_387_n N_B_c_579_n 6.16253e-19
cc_282 N_A_c_379_n B 7.07944e-19
cc_283 N_A_c_387_n B 5.00495e-19
cc_284 N_A_c_379_n N_B_c_615_n 2.41829e-19
cc_285 N_A_c_401_n N_B_c_583_n 8.44727e-19
cc_286 N_A_c_434_p N_B_c_583_n 4.84491e-19
cc_287 N_A_c_378_n N_B_c_580_n 2.87365e-19
cc_288 N_A_c_387_n N_B_c_580_n 6.85754e-19
cc_289 N_A_c_379_n N_B_c_620_n 3.8563e-19
cc_290 N_A_XI3.X0_PGD N_B_c_621_n 0.00133285f
cc_291 N_A_c_401_n N_B_c_621_n 4.67029e-19
cc_292 N_A_c_434_p N_B_c_621_n 0.0014909f
cc_293 N_A_c_387_n N_B_c_581_n 0.00225059f
cc_294 N_A_c_396_n N_B_c_581_n 8.88958e-19
cc_295 N_A_c_379_n N_B_c_602_n 0.00244205f
cc_296 N_A_c_396_n N_Z_XI2.X0_D 6.94686e-19
cc_297 N_A_XI3.X0_PGD N_Z_c_669_n 6.30408e-19
cc_298 N_A_c_387_n N_Z_c_669_n 0.00124827f
cc_299 N_A_c_396_n N_Z_c_669_n 0.00121415f
cc_300 N_BI_XI2.X0_CG N_AI_XI2.X0_PGD 8.63152e-19
cc_301 N_BI_c_486_n N_AI_XI2.X0_PGD 0.00133285f
cc_302 N_BI_c_464_n N_AI_c_529_n 3.64122e-19
cc_303 N_BI_c_464_n N_B_c_579_n 0.00139574f
cc_304 N_BI_c_464_n N_B_c_615_n 6.02887e-19
cc_305 N_BI_c_479_n N_B_c_615_n 3.05615e-19
cc_306 N_BI_c_478_n N_B_c_583_n 0.00178808f
cc_307 N_BI_c_467_n N_B_c_583_n 0.00156529f
cc_308 N_BI_c_464_n N_B_c_620_n 4.56568e-19
cc_309 N_BI_c_486_n N_B_c_620_n 0.00266354f
cc_310 N_BI_c_487_n N_B_c_620_n 7.16621e-19
cc_311 N_BI_c_478_n N_B_c_621_n 4.56568e-19
cc_312 N_BI_c_486_n N_B_c_621_n 6.17967e-19
cc_313 N_BI_c_487_n N_B_c_621_n 0.00243716f
cc_314 N_BI_c_464_n N_B_c_581_n 0.00427216f
cc_315 N_BI_c_464_n N_B_c_603_n 3.15526e-19
cc_316 N_BI_c_467_n N_B_c_603_n 0.00129112f
cc_317 N_BI_c_506_p N_B_c_603_n 0.0034245f
cc_318 N_BI_c_464_n N_B_c_585_n 4.99817e-19
cc_319 N_BI_c_467_n N_B_c_585_n 7.12768e-19
cc_320 N_BI_c_479_n N_B_c_585_n 7.15853e-19
cc_321 N_BI_c_506_p N_B_c_645_n 0.00229162f
cc_322 N_BI_c_464_n N_B_c_586_n 0.00139788f
cc_323 N_BI_c_467_n N_B_c_586_n 8.65145e-19
cc_324 N_BI_c_464_n N_Z_c_669_n 0.00138937f
cc_325 N_BI_c_478_n N_Z_c_669_n 0.00157561f
cc_326 N_BI_c_486_n N_Z_c_669_n 8.66889e-19
cc_327 N_BI_c_467_n N_Z_c_669_n 0.00100271f
cc_328 N_BI_c_506_p N_Z_c_669_n 0.00210866f
cc_329 N_BI_c_479_n N_Z_c_669_n 9.67357e-19
cc_330 N_AI_XI2.X0_PGD N_B_c_648_n 8.79767e-19
cc_331 N_AI_c_527_n N_B_c_648_n 0.00234569f
cc_332 N_AI_c_537_n N_B_c_615_n 5.49665e-19
cc_333 N_AI_c_527_n N_B_c_615_n 4.745e-19
cc_334 N_AI_XI2.X0_PGD N_B_c_620_n 0.00133285f
cc_335 N_AI_c_566_p N_B_c_620_n 7.60534e-19
cc_336 N_AI_c_537_n N_B_c_620_n 4.46045e-19
cc_337 N_AI_c_527_n N_B_c_620_n 0.00166302f
cc_338 N_AI_c_528_n N_B_c_581_n 0.00120142f
cc_339 N_AI_c_529_n N_B_c_581_n 3.28172e-19
cc_340 N_AI_c_529_n N_B_c_602_n 2.8335e-19
cc_341 N_AI_c_537_n N_B_c_603_n 4.27113e-19
cc_342 N_AI_XI2.X0_PGD N_Z_c_669_n 3.26804e-19
cc_343 N_B_c_615_n N_Z_c_669_n 0.0013937f
cc_344 N_B_c_583_n N_Z_c_669_n 0.00139745f
cc_345 N_B_c_620_n N_Z_c_669_n 8.66889e-19
cc_346 N_B_c_621_n N_Z_c_669_n 8.66889e-19
cc_347 N_B_c_603_n N_Z_c_669_n 4.72173e-19
*
.ends
*
*
.subckt XOR3_HPNW4 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XOR3_N1
.ends
