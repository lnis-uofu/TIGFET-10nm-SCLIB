* sclib_tigfet10_hpnw12_tt_0p70v_25c.sp
.subckt TIGFET_HPNW12 D PGD CG PGS S
xgate (D PGD CG PGS S) TIGFET nw=12
.ends
*
* File: G3_AND2_N3.pex.netlist
* Created: Tue Mar  1 10:56:10 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_AND2_N3_VSS 2 4 6 8 10 12 14 16 30 31 50 62 67 70 75 80 85 94 99
+ 108 109 113 114 119 125 127 132 133 134 136 Vss
c67 134 Vss 3.75522e-19
c68 133 Vss 3.62111e-19
c69 132 Vss 0.004799f
c70 127 Vss 0.00257088f
c71 125 Vss 0.00552282f
c72 119 Vss 0.00412002f
c73 114 Vss 8.41284e-19
c74 113 Vss 0.00175777f
c75 109 Vss 7.31223e-19
c76 108 Vss 0.00590165f
c77 99 Vss 0.00416928f
c78 94 Vss 0.00536429f
c79 85 Vss 7.10513e-22
c80 80 Vss 4.8997e-19
c81 75 Vss 0.00125499f
c82 70 Vss 0.00121927f
c83 67 Vss 0.0100822f
c84 62 Vss 0.00955849f
c85 58 Vss 0.0299311f
c86 57 Vss 0.0299311f
c87 51 Vss 0.0357161f
c88 50 Vss 0.0994129f
c89 42 Vss 0.107716f
c90 37 Vss 0.0688416f
c91 31 Vss 0.0350852f
c92 30 Vss 0.0646396f
c93 14 Vss 0.188821f
c94 12 Vss 0.189513f
c95 10 Vss 0.189371f
c96 8 Vss 0.190733f
c97 6 Vss 0.189919f
c98 4 Vss 0.190281f
c99 2 Vss 1.99696e-19
r100 132 136 0.326018
r101 131 132 5.50157
r102 127 131 0.655813
r103 126 134 0.494161
r104 125 136 0.326018
r105 125 126 10.1279
r106 121 134 0.128424
r107 120 133 0.494161
r108 119 134 0.494161
r109 119 120 10.378
r110 115 133 0.128424
r111 113 133 0.494161
r112 113 114 4.33457
r113 108 114 0.652036
r114 107 109 0.655813
r115 107 108 19.0471
r116 85 127 1.82344
r117 80 99 1.16709
r118 80 121 2.16729
r119 75 94 1.16709
r120 75 115 2.16729
r121 70 109 1.82344
r122 67 85 1.16709
r123 62 70 1.16709
r124 53 99 0.0476429
r125 51 53 1.45875
r126 50 54 0.652036
r127 50 53 1.45875
r128 47 51 0.652036
r129 43 58 0.494161
r130 42 44 0.652036
r131 42 43 2.9175
r132 39 58 0.128424
r133 38 57 0.494161
r134 37 58 0.494161
r135 37 38 2.8008
r136 34 57 0.128424
r137 33 94 0.0476429
r138 31 33 1.4004
r139 30 57 0.494161
r140 30 33 1.5171
r141 27 31 0.652036
r142 16 67 0.123773
r143 14 47 5.1348
r144 12 54 5.1348
r145 10 44 5.1348
r146 8 39 5.1348
r147 6 27 5.1348
r148 4 34 5.1348
r149 2 62 0.123773
.ends

.subckt PM_G3_AND2_N3_VDD 2 4 6 8 10 12 25 27 33 43 48 51 53 54 58 60 64 68 70
+ 74 76 78 79 85 94 Vss
c86 94 Vss 0.00463585f
c87 85 Vss 0.00402796f
c88 79 Vss 4.43941e-19
c89 76 Vss 4.52364e-19
c90 74 Vss 7.90245e-19
c91 70 Vss 0.00408718f
c92 68 Vss 0.00117255f
c93 64 Vss 0.00432275f
c94 60 Vss 0.00739867f
c95 58 Vss 0.00173558f
c96 55 Vss 0.00171371f
c97 54 Vss 0.0100369f
c98 53 Vss 0.00360598f
c99 51 Vss 0.00814794f
c100 48 Vss 0.00687623f
c101 43 Vss 0.00811526f
c102 33 Vss 0.0357902f
c103 32 Vss 0.102427f
c104 27 Vss 0.170038f
c105 25 Vss 0.0352365f
c106 12 Vss 0.190935f
c107 10 Vss 0.189512f
c108 8 Vss 0.00143493f
c109 2 Vss 0.221827f
r110 74 94 1.16709
r111 72 74 2.16729
r112 71 79 0.494161
r113 70 72 0.652036
r114 70 71 7.46046
r115 66 79 0.128424
r116 66 68 6.16843
r117 64 85 1.16709
r118 62 64 6.08507
r119 61 78 0.326018
r120 60 79 0.494161
r121 60 61 13.0037
r122 56 76 0.0828784
r123 56 58 1.82344
r124 54 62 0.652036
r125 54 55 10.0862
r126 53 78 0.326018
r127 52 76 0.551426
r128 52 53 5.50157
r129 51 76 0.551426
r130 50 55 0.652036
r131 50 51 15.046
r132 48 68 1.16709
r133 43 58 1.16709
r134 35 94 0.0476429
r135 33 35 1.45875
r136 32 36 0.652036
r137 32 35 1.45875
r138 29 33 0.652036
r139 27 85 0.428786
r140 25 27 5.3682
r141 22 25 0.652036
r142 12 36 5.1348
r143 10 29 5.1348
r144 8 48 0.123773
r145 6 48 0.123773
r146 4 43 0.123773
r147 2 22 6.3018
.ends

.subckt PM_G3_AND2_N3_A 1 2 9 20 23 28 33 Vss
c24 33 Vss 0.00369912f
c25 28 Vss 0.00225353f
c26 20 Vss 0.00104617f
c27 12 Vss 0.166756f
c28 1 Vss 0.171396f
r29 25 33 1.16709
r30 23 25 2.66743
r31 20 28 1.16709
r32 20 23 2.70911
r33 12 33 0.50025
r34 9 28 0.50025
r35 2 12 4.37625
r36 1 9 4.60965
.ends

.subckt PM_G3_AND2_N3_NET1 2 4 6 7 8 23 26 38 42 48 52 54 58 71 Vss
c52 71 Vss 0.00600165f
c53 60 Vss 2.11292e-19
c54 58 Vss 0.0011885f
c55 54 Vss 0.00636228f
c56 52 Vss 6.44544e-19
c57 48 Vss 8.20028e-19
c58 42 Vss 0.00560082f
c59 38 Vss 0.00901424f
c60 26 Vss 8.44333e-20
c61 23 Vss 0.229828f
c62 19 Vss 0.18045f
c63 17 Vss 0.0247918f
c64 8 Vss 0.193588f
c65 6 Vss 0.00143493f
r66 58 71 1.16709
r67 56 58 2.16729
r68 55 60 0.128424
r69 54 56 0.652036
r70 54 55 7.46046
r71 52 68 1.16709
r72 50 60 0.494161
r73 50 52 6.29346
r74 46 60 0.494161
r75 46 48 6.21011
r76 42 68 0.15
r77 38 48 1.16709
r78 26 71 0.0476429
r79 24 26 0.326018
r80 24 26 0.1167
r81 23 27 0.652036
r82 23 26 6.7686
r83 19 71 0.357321
r84 17 26 0.326018
r85 17 19 0.40845
r86 8 27 5.1348
r87 7 19 4.72635
r88 6 42 0.123773
r89 4 42 0.123773
r90 2 38 0.123773
.ends

.subckt PM_G3_AND2_N3_B 2 3 9 10 13 19 22 Vss
c26 19 Vss 2.97116e-19
c27 13 Vss 0.236449f
c28 10 Vss 0.0348969f
c29 9 Vss 0.287374f
c30 2 Vss 0.332764f
r31 19 22 0.0416786
r32 13 19 1.16709
r33 11 13 2.15895
r34 9 11 0.652036
r35 9 10 8.92755
r36 6 10 0.652036
r37 3 13 5.6016
r38 2 6 10.0362
.ends

.subckt PM_G3_AND2_N3_Z 2 4 13 16 Vss
c13 13 Vss 0.00498872f
c14 4 Vss 0.00143493f
r15 16 19 0.0416786
r16 13 19 1.16709
r17 4 13 0.123773
r18 2 13 0.123773
.ends

.subckt G3_AND2_N3  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI13.X0 N_NET1_XI13.X0_D N_VDD_XI13.X0_PGD N_A_XI13.X0_CG N_B_XI13.X0_PGS
+ N_VSS_XI13.X0_S TIGFET_HPNW12
XI15.X0 N_NET1_XI15.X0_D N_VSS_XI15.X0_PGD N_A_XI15.X0_CG N_VSS_XI15.X0_PGS
+ N_VDD_XI15.X0_S TIGFET_HPNW12
XI14.X0 N_NET1_XI14.X0_D N_VSS_XI14.X0_PGD N_B_XI14.X0_CG N_VSS_XI14.X0_PGS
+ N_VDD_XI14.X0_S TIGFET_HPNW12
XI12.X0 N_Z_XI12.X0_D N_VSS_XI12.X0_PGD N_NET1_XI12.X0_CG N_VSS_XI12.X0_PGS
+ N_VDD_XI12.X0_S TIGFET_HPNW12
XI11.X0 N_Z_XI11.X0_D N_VDD_XI11.X0_PGD N_NET1_XI11.X0_CG N_VDD_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW12
*
x_PM_G3_AND2_N3_VSS N_VSS_XI13.X0_S N_VSS_XI15.X0_PGD N_VSS_XI15.X0_PGS
+ N_VSS_XI14.X0_PGD N_VSS_XI14.X0_PGS N_VSS_XI12.X0_PGD N_VSS_XI12.X0_PGS
+ N_VSS_XI11.X0_S N_VSS_c_14_p N_VSS_c_15_p N_VSS_c_2_p N_VSS_c_3_p N_VSS_c_62_p
+ N_VSS_c_4_p N_VSS_c_8_p N_VSS_c_24_p N_VSS_c_63_p N_VSS_c_9_p N_VSS_c_26_p
+ N_VSS_c_5_p N_VSS_c_6_p N_VSS_c_18_p N_VSS_c_11_p N_VSS_c_19_p N_VSS_c_33_p
+ N_VSS_c_67_p N_VSS_c_28_p N_VSS_c_20_p N_VSS_c_34_p VSS Vss PM_G3_AND2_N3_VSS
x_PM_G3_AND2_N3_VDD N_VDD_XI13.X0_PGD N_VDD_XI15.X0_S N_VDD_XI14.X0_S
+ N_VDD_XI12.X0_S N_VDD_XI11.X0_PGD N_VDD_XI11.X0_PGS N_VDD_c_146_p
+ N_VDD_c_128_p N_VDD_c_69_n N_VDD_c_122_p N_VDD_c_123_p N_VDD_c_70_n
+ N_VDD_c_74_n N_VDD_c_79_n N_VDD_c_80_n N_VDD_c_81_n N_VDD_c_121_p N_VDD_c_88_n
+ N_VDD_c_96_n N_VDD_c_102_n N_VDD_c_105_n VDD N_VDD_c_106_n N_VDD_c_117_p
+ N_VDD_c_107_n Vss PM_G3_AND2_N3_VDD
x_PM_G3_AND2_N3_A N_A_XI13.X0_CG N_A_XI15.X0_CG N_A_c_160_n N_A_c_154_n A
+ N_A_c_163_n N_A_c_156_n Vss PM_G3_AND2_N3_A
x_PM_G3_AND2_N3_NET1 N_NET1_XI13.X0_D N_NET1_XI15.X0_D N_NET1_XI14.X0_D
+ N_NET1_XI12.X0_CG N_NET1_XI11.X0_CG N_NET1_c_178_n N_NET1_c_179_n
+ N_NET1_c_180_n N_NET1_c_194_n N_NET1_c_182_n N_NET1_c_185_n N_NET1_c_186_n
+ N_NET1_c_188_n N_NET1_c_190_n Vss PM_G3_AND2_N3_NET1
x_PM_G3_AND2_N3_B N_B_XI13.X0_PGS N_B_XI14.X0_CG N_B_c_230_n N_B_c_232_n
+ N_B_c_237_n N_B_c_252_n B Vss PM_G3_AND2_N3_B
x_PM_G3_AND2_N3_Z N_Z_XI12.X0_D N_Z_XI11.X0_D N_Z_c_256_n Z Vss PM_G3_AND2_N3_Z
cc_1 N_VSS_XI12.X0_PGD N_VDD_XI11.X0_PGD 0.00195824f
cc_2 N_VSS_c_2_p N_VDD_c_69_n 0.00195824f
cc_3 N_VSS_c_3_p N_VDD_c_70_n 9.5668e-19
cc_4 N_VSS_c_4_p N_VDD_c_70_n 0.00165395f
cc_5 N_VSS_c_5_p N_VDD_c_70_n 0.00795264f
cc_6 N_VSS_c_6_p N_VDD_c_70_n 0.00190019f
cc_7 N_VSS_XI15.X0_PGS N_VDD_c_74_n 3.39564e-19
cc_8 N_VSS_c_8_p N_VDD_c_74_n 4.42007e-19
cc_9 N_VSS_c_9_p N_VDD_c_74_n 3.70842e-19
cc_10 N_VSS_c_5_p N_VDD_c_74_n 0.00357958f
cc_11 N_VSS_c_11_p N_VDD_c_74_n 0.00107567f
cc_12 N_VSS_c_4_p N_VDD_c_79_n 0.00237483f
cc_13 N_VSS_c_4_p N_VDD_c_80_n 3.67743e-19
cc_14 N_VSS_c_14_p N_VDD_c_81_n 0.00161328f
cc_15 N_VSS_c_15_p N_VDD_c_81_n 3.76573e-19
cc_16 N_VSS_c_8_p N_VDD_c_81_n 0.00161703f
cc_17 N_VSS_c_9_p N_VDD_c_81_n 2.26455e-19
cc_18 N_VSS_c_18_p N_VDD_c_81_n 0.00349492f
cc_19 N_VSS_c_19_p N_VDD_c_81_n 0.00593063f
cc_20 N_VSS_c_20_p N_VDD_c_81_n 7.61747e-19
cc_21 N_VSS_XI14.X0_PGS N_VDD_c_88_n 2.0368e-19
cc_22 N_VSS_XI12.X0_PGS N_VDD_c_88_n 2.24983e-19
cc_23 N_VSS_c_8_p N_VDD_c_88_n 6.58919e-19
cc_24 N_VSS_c_24_p N_VDD_c_88_n 0.0018079f
cc_25 N_VSS_c_9_p N_VDD_c_88_n 2.56577e-19
cc_26 N_VSS_c_26_p N_VDD_c_88_n 9.55109e-19
cc_27 N_VSS_c_5_p N_VDD_c_88_n 4.30333e-19
cc_28 N_VSS_c_28_p N_VDD_c_88_n 2.91233e-19
cc_29 N_VSS_c_2_p N_VDD_c_96_n 5.15102e-19
cc_30 N_VSS_c_24_p N_VDD_c_96_n 0.00161703f
cc_31 N_VSS_c_26_p N_VDD_c_96_n 2.26455e-19
cc_32 N_VSS_c_19_p N_VDD_c_96_n 0.00133474f
cc_33 N_VSS_c_33_p N_VDD_c_96_n 0.00600556f
cc_34 N_VSS_c_34_p N_VDD_c_96_n 7.74609e-19
cc_35 N_VSS_c_24_p N_VDD_c_102_n 8.50587e-19
cc_36 N_VSS_c_26_p N_VDD_c_102_n 3.82294e-19
cc_37 N_VSS_c_28_p N_VDD_c_102_n 3.85245e-19
cc_38 N_VSS_c_5_p N_VDD_c_105_n 0.00100712f
cc_39 N_VSS_c_19_p N_VDD_c_106_n 9.82771e-19
cc_40 N_VSS_c_24_p N_VDD_c_107_n 3.48267e-19
cc_41 N_VSS_c_26_p N_VDD_c_107_n 6.46219e-19
cc_42 N_VSS_c_9_p N_A_c_154_n 2.354e-19
cc_43 N_VSS_c_5_p N_A_c_154_n 0.00149458f
cc_44 N_VSS_c_8_p N_A_c_156_n 2.15082e-19
cc_45 N_VSS_c_9_p N_A_c_156_n 4.9359e-19
cc_46 N_VSS_XI12.X0_PGD N_NET1_c_178_n 4.31283e-19
cc_47 N_VSS_c_26_p N_NET1_c_179_n 5.28949e-19
cc_48 N_VSS_c_3_p N_NET1_c_180_n 3.43419e-19
cc_49 N_VSS_c_4_p N_NET1_c_180_n 3.48267e-19
cc_50 N_VSS_c_3_p N_NET1_c_182_n 3.48267e-19
cc_51 N_VSS_c_4_p N_NET1_c_182_n 8.50248e-19
cc_52 N_VSS_c_5_p N_NET1_c_182_n 8.95101e-19
cc_53 N_VSS_c_19_p N_NET1_c_185_n 2.278e-19
cc_54 N_VSS_XI14.X0_PGS N_NET1_c_186_n 2.25423e-19
cc_55 N_VSS_c_19_p N_NET1_c_186_n 4.57847e-19
cc_56 N_VSS_c_24_p N_NET1_c_188_n 2.00623e-19
cc_57 N_VSS_c_26_p N_NET1_c_188_n 2.28697e-19
cc_58 N_VSS_c_24_p N_NET1_c_190_n 2.15082e-19
cc_59 N_VSS_XI15.X0_PGD N_B_c_230_n 8.16475e-19
cc_60 N_VSS_XI14.X0_PGD N_B_c_230_n 8.16475e-19
cc_61 N_VSS_XI15.X0_PGS N_B_c_232_n 0.00101175f
cc_62 N_VSS_c_62_p N_Z_c_256_n 3.43419e-19
cc_63 N_VSS_c_63_p N_Z_c_256_n 3.48267e-19
cc_64 N_VSS_c_62_p Z 3.48267e-19
cc_65 N_VSS_c_63_p Z 4.99861e-19
cc_66 N_VSS_c_33_p Z 2.23989e-19
cc_67 N_VSS_c_67_p Z 2.7826e-19
cc_68 N_VDD_XI13.X0_PGD N_A_XI13.X0_CG 4.85665e-19
cc_69 N_VDD_c_79_n N_A_XI13.X0_CG 3.10124e-19
cc_70 N_VDD_c_79_n N_A_c_160_n 2.67445e-19
cc_71 N_VDD_c_70_n N_A_c_154_n 0.0028804f
cc_72 N_VDD_c_79_n N_A_c_154_n 4.70376e-19
cc_73 N_VDD_XI13.X0_PGD N_A_c_163_n 4.86892e-19
cc_74 N_VDD_c_70_n N_A_c_163_n 3.66936e-19
cc_75 N_VDD_c_79_n N_A_c_163_n 2.64879e-19
cc_76 N_VDD_c_117_p N_A_c_163_n 5.21476e-19
cc_77 N_VDD_c_70_n N_A_c_156_n 5.07754e-19
cc_78 N_VDD_XI11.X0_PGD N_NET1_c_178_n 4.31283e-19
cc_79 N_VDD_c_79_n N_NET1_c_180_n 0.0011619f
cc_80 N_VDD_c_121_p N_NET1_c_180_n 8.835e-19
cc_81 N_VDD_c_122_p N_NET1_c_194_n 3.43419e-19
cc_82 N_VDD_c_123_p N_NET1_c_194_n 3.43419e-19
cc_83 N_VDD_c_80_n N_NET1_c_194_n 3.72199e-19
cc_84 N_VDD_c_81_n N_NET1_c_194_n 2.82909e-19
cc_85 N_VDD_c_88_n N_NET1_c_194_n 3.48267e-19
cc_86 N_VDD_XI13.X0_PGD N_NET1_c_182_n 3.17068e-19
cc_87 N_VDD_c_128_p N_NET1_c_182_n 8.01918e-19
cc_88 N_VDD_c_70_n N_NET1_c_182_n 0.00133415f
cc_89 N_VDD_c_79_n N_NET1_c_182_n 0.00168724f
cc_90 N_VDD_c_121_p N_NET1_c_182_n 0.00619213f
cc_91 N_VDD_c_117_p N_NET1_c_182_n 9.07013e-19
cc_92 N_VDD_c_122_p N_NET1_c_185_n 3.48267e-19
cc_93 N_VDD_c_123_p N_NET1_c_185_n 3.48267e-19
cc_94 N_VDD_c_80_n N_NET1_c_185_n 8.08807e-19
cc_95 N_VDD_c_81_n N_NET1_c_185_n 3.96039e-19
cc_96 N_VDD_c_88_n N_NET1_c_185_n 7.82265e-19
cc_97 N_VDD_c_128_p N_NET1_c_186_n 3.89384e-19
cc_98 N_VDD_c_123_p N_NET1_c_186_n 2.74986e-19
cc_99 N_VDD_c_121_p N_NET1_c_186_n 0.00138769f
cc_100 N_VDD_c_88_n N_NET1_c_186_n 5.47694e-19
cc_101 N_VDD_c_117_p N_NET1_c_186_n 8.66889e-19
cc_102 N_VDD_XI13.X0_PGD N_B_XI13.X0_PGS 0.00331493f
cc_103 N_VDD_c_70_n N_B_XI13.X0_PGS 7.63549e-19
cc_104 N_VDD_c_79_n N_B_XI13.X0_PGS 6.44483e-19
cc_105 N_VDD_c_146_p N_B_c_230_n 0.00792574f
cc_106 N_VDD_c_117_p N_B_c_237_n 0.0014275f
cc_107 N_VDD_c_123_p N_Z_c_256_n 3.43419e-19
cc_108 N_VDD_c_88_n N_Z_c_256_n 3.48267e-19
cc_109 N_VDD_c_96_n N_Z_c_256_n 2.74986e-19
cc_110 N_VDD_c_123_p Z 3.48267e-19
cc_111 N_VDD_c_88_n Z 7.09569e-19
cc_112 N_VDD_c_96_n Z 3.66281e-19
cc_113 N_A_c_154_n N_NET1_c_182_n 0.0080879f
cc_114 N_A_c_163_n N_NET1_c_182_n 8.85473e-19
cc_115 N_A_c_156_n N_NET1_c_185_n 9.58642e-19
cc_116 N_A_XI13.X0_CG N_B_XI13.X0_PGS 4.84447e-19
cc_117 N_A_c_154_n N_B_XI13.X0_PGS 3.59952e-19
cc_118 N_A_c_163_n N_B_XI13.X0_PGS 5.64689e-19
cc_119 N_A_c_154_n N_B_c_230_n 2.067e-19
cc_120 N_A_c_163_n N_B_c_230_n 6.90429e-19
cc_121 N_A_c_156_n N_B_c_230_n 0.0015879f
cc_122 N_A_c_156_n N_B_c_237_n 9.27569e-19
cc_123 N_NET1_c_194_n N_B_c_230_n 3.4562e-19
cc_124 N_NET1_c_185_n N_B_c_230_n 2.39796e-19
cc_125 N_NET1_c_186_n N_B_c_230_n 4.12724e-19
cc_126 N_NET1_c_185_n N_B_c_237_n 0.00116203f
cc_127 N_NET1_c_186_n N_B_c_237_n 0.00112058f
cc_128 N_NET1_c_188_n N_B_c_237_n 3.86148e-19
cc_129 N_NET1_c_190_n N_B_c_237_n 0.00196155f
cc_130 N_NET1_c_185_n N_B_c_252_n 0.00147455f
cc_131 N_NET1_c_186_n N_B_c_252_n 0.00146537f
cc_132 N_NET1_c_188_n N_B_c_252_n 5.75904e-19
cc_133 N_NET1_c_190_n N_B_c_252_n 3.48267e-19
cc_134 N_NET1_c_178_n N_Z_c_256_n 7.69306e-19
*
.ends
*
*
.subckt AND2_HPNW12 A B Y VDD VSS
xgate (VSS VDD A B Y) G3_AND2_N3
.ends
*
* File: G2_AOI21_N3.pex.netlist
* Created: Mon Apr 11 18:50:47 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_AOI21_N3_VSS 2 4 6 8 19 30 35 38 43 48 57 66 67 69 77 78 79 84 86
+ 88 89 Vss
c48 89 Vss 4.28045e-19
c49 86 Vss 0.00576702f
c50 84 Vss 0.00198426f
c51 79 Vss 0.00132518f
c52 78 Vss 4.66086e-19
c53 77 Vss 0.00250771f
c54 69 Vss 0.00104615f
c55 67 Vss 0.0101744f
c56 66 Vss 0.00354326f
c57 65 Vss 0.00133883f
c58 57 Vss 0.00699915f
c59 48 Vss 2.01624e-19
c60 43 Vss 0.00190058f
c61 38 Vss 0.00140655f
c62 35 Vss 0.00813966f
c63 30 Vss 0.0101549f
c64 25 Vss 0.0829032f
c65 19 Vss 0.0350566f
c66 18 Vss 0.0688416f
c67 8 Vss 0.190897f
c68 4 Vss 0.189497f
r69 85 89 0.551426
r70 85 86 18.3386
r71 84 89 0.551426
r72 83 84 5.50157
r73 79 89 0.0828784
r74 77 86 0.652036
r75 77 78 4.33457
r76 73 78 0.652036
r77 68 88 0.326149
r78 67 83 0.652298
r79 67 68 15.1308
r80 66 69 0.655813
r81 65 88 0.326149
r82 65 66 5.50157
r83 48 79 1.82344
r84 43 57 1.16709
r85 43 73 2.16729
r86 38 69 1.82344
r87 35 48 1.16709
r88 30 38 1.16709
r89 25 57 0.0476429
r90 23 25 2.04225
r91 20 23 0.0685365
r92 18 23 0.5835
r93 18 19 2.8008
r94 15 19 0.652036
r95 8 20 5.1348
r96 6 35 0.123773
r97 4 15 5.1348
r98 2 30 0.123773
.ends

.subckt PM_G2_AOI21_N3_VDD 2 4 6 8 10 29 37 42 45 46 48 50 54 56 57 58 63 65 66
+ 68 74 Vss
c56 74 Vss 0.004704f
c57 66 Vss 4.52364e-19
c58 65 Vss 0.00371658f
c59 63 Vss 0.0104139f
c60 58 Vss 0.0017471f
c61 57 Vss 6.04409e-19
c62 56 Vss 0.00309603f
c63 54 Vss 0.00137895f
c64 51 Vss 0.00173381f
c65 50 Vss 0.0117653f
c66 48 Vss 0.00158874f
c67 46 Vss 0.00143356f
c68 45 Vss 0.00419705f
c69 42 Vss 0.0082636f
c70 37 Vss 0.010107f
c71 33 Vss 0.0307825f
c72 29 Vss 8.92604e-20
c73 26 Vss 0.101624f
c74 22 Vss 0.0359157f
c75 21 Vss 0.0712517f
c76 8 Vss 0.189919f
c77 6 Vss 0.190671f
c78 2 Vss 0.189552f
r79 65 68 0.326018
r80 64 66 0.551426
r81 64 65 5.50157
r82 63 66 0.551426
r83 62 63 18.3386
r84 58 66 0.0828784
r85 58 60 1.82344
r86 56 62 0.652036
r87 56 57 4.37625
r88 54 74 1.16709
r89 52 57 0.652036
r90 52 54 2.16729
r91 50 68 0.326018
r92 50 51 15.6711
r93 46 48 1.82344
r94 45 51 0.652036
r95 44 46 0.655813
r96 44 45 5.50157
r97 42 60 1.16709
r98 37 48 1.16709
r99 29 74 0.0476429
r100 27 33 0.494161
r101 27 29 1.45875
r102 26 30 0.652036
r103 26 29 1.45875
r104 23 33 0.128424
r105 21 33 0.494161
r106 21 22 2.8008
r107 18 22 0.652036
r108 10 42 0.123773
r109 8 30 5.1348
r110 6 23 5.1348
r111 4 37 0.123773
r112 2 18 5.1348
.ends

.subckt PM_G2_AOI21_N3_B 2 4 20 23 26 29 Vss
c18 29 Vss 0.00496711f
c19 23 Vss 4.14813e-19
c20 20 Vss 0.0923936f
c21 16 Vss 0.0610957f
c22 4 Vss 0.211686f
c23 2 Vss 0.427124f
r24 23 29 1.16709
r25 23 26 0.125036
r26 18 20 2.04225
r27 16 29 0.197068
r28 13 16 1.2837
r29 10 20 0.0685365
r30 8 18 0.0685365
r31 7 13 0.0685365
r32 4 10 5.6016
r33 2 8 11.2032
r34 2 7 5.1348
.ends

.subckt PM_G2_AOI21_N3_C 2 4 6 17 24 28 31 36 39 43 56 Vss
c47 56 Vss 0.00111429f
c48 43 Vss 0.0052438f
c49 39 Vss 0.00260114f
c50 36 Vss 3.26162e-19
c51 31 Vss 0.00720813f
c52 28 Vss 0.0949366f
c53 24 Vss 0.084323f
c54 17 Vss 4.93054e-19
c55 6 Vss 0.286419f
c56 4 Vss 0.25621f
c57 2 Vss 0.189817f
r58 52 56 0.652036
r59 39 56 5.16814
r60 36 39 0.0833571
r61 31 43 1.16709
r62 31 52 12.2535
r63 26 28 2.04225
r64 24 43 0.0476429
r65 21 24 1.92555
r66 18 28 0.0685365
r67 17 39 1.16709
r68 13 26 0.0685365
r69 13 17 2.8008
r70 10 21 0.0685365
r71 6 18 8.4024
r72 4 17 5.6016
r73 2 10 5.1348
.ends

.subckt PM_G2_AOI21_N3_Z 2 4 6 8 23 27 30 33 Vss
c33 30 Vss 0.00262006f
c34 27 Vss 0.00473513f
c35 23 Vss 0.00644988f
c36 8 Vss 0.00143493f
c37 6 Vss 0.00143493f
r38 33 35 7.5855
r39 30 33 5.2515
r40 27 35 1.16709
r41 23 30 1.16709
r42 8 27 0.123773
r43 6 23 0.123773
r44 4 27 0.123773
r45 2 23 0.123773
.ends

.subckt PM_G2_AOI21_N3_A 2 4 10 11 13 14 15 20 24 29 32 Vss
c32 32 Vss 9.42706e-19
c33 29 Vss 5.87748e-19
c34 24 Vss 1.66175e-19
c35 20 Vss 0.191363f
c36 18 Vss 0.0247918f
c37 15 Vss 0.0322409f
c38 14 Vss 0.0740343f
c39 13 Vss 0.0312529f
c40 11 Vss 0.0324985f
c41 10 Vss 0.122088f
c42 2 Vss 0.292885f
r43 26 32 1.16709
r44 26 29 0.0729375
r45 24 32 0.262036
r46 20 32 0.238214
r47 18 24 0.326018
r48 18 20 0.64185
r49 15 24 2.50905
r50 14 24 0.326018
r51 14 24 0.1167
r52 13 15 0.652036
r53 12 13 1.22535
r54 10 12 0.652036
r55 10 11 3.09255
r56 7 11 0.652036
r57 4 20 5.0181
r58 2 7 8.7525
.ends

.subckt G2_AOI21_N3  VSS VDD B C Z A
*
* A	A
* Z	Z
* C	C
* B	B
* VDD	VDD
* VSS	VSS
XI18.X0 N_Z_XI18.X0_D N_VDD_XI18.X0_PGD N_A_XI18.X0_CG N_B_XI18.X0_PGS
+ N_VSS_XI18.X0_S TIGFET_HPNW12
XI16.X0 N_Z_XI16.X0_D N_VSS_XI16.X0_PGD N_B_XI16.X0_CG N_C_XI16.X0_PGS
+ N_VDD_XI16.X0_S TIGFET_HPNW12
XI19.X0 N_Z_XI19.X0_D N_VDD_XI19.X0_PGD N_C_XI19.X0_CG N_VDD_XI19.X0_PGS
+ N_VSS_XI19.X0_S TIGFET_HPNW12
XI17.X0 N_Z_XI17.X0_D N_VSS_XI17.X0_PGD N_A_XI17.X0_CG N_C_XI17.X0_PGS
+ N_VDD_XI17.X0_S TIGFET_HPNW12
*
x_PM_G2_AOI21_N3_VSS N_VSS_XI18.X0_S N_VSS_XI16.X0_PGD N_VSS_XI19.X0_S
+ N_VSS_XI17.X0_PGD N_VSS_c_3_p N_VSS_c_34_p N_VSS_c_8_p N_VSS_c_2_p N_VSS_c_4_p
+ N_VSS_c_9_p N_VSS_c_5_p N_VSS_c_21_p N_VSS_c_10_p N_VSS_c_1_p N_VSS_c_6_p
+ N_VSS_c_7_p N_VSS_c_12_p N_VSS_c_14_p N_VSS_c_15_p VSS N_VSS_c_16_p Vss
+ PM_G2_AOI21_N3_VSS
x_PM_G2_AOI21_N3_VDD N_VDD_XI18.X0_PGD N_VDD_XI16.X0_S N_VDD_XI19.X0_PGD
+ N_VDD_XI19.X0_PGS N_VDD_XI17.X0_S N_VDD_c_76_p N_VDD_c_90_p N_VDD_c_91_p
+ N_VDD_c_75_p N_VDD_c_49_n N_VDD_c_50_n N_VDD_c_51_n N_VDD_c_70_p N_VDD_c_56_n
+ N_VDD_c_59_n N_VDD_c_60_n N_VDD_c_61_n N_VDD_c_65_n N_VDD_c_68_n VDD
+ N_VDD_c_71_p Vss PM_G2_AOI21_N3_VDD
x_PM_G2_AOI21_N3_B N_B_XI18.X0_PGS N_B_XI16.X0_CG N_B_c_113_p N_B_c_105_n B
+ N_B_c_110_n Vss PM_G2_AOI21_N3_B
x_PM_G2_AOI21_N3_C N_C_XI16.X0_PGS N_C_XI19.X0_CG N_C_XI17.X0_PGS N_C_c_135_n
+ N_C_c_137_n N_C_c_138_n N_C_c_124_n C N_C_c_127_n N_C_c_128_n N_C_c_132_n Vss
+ PM_G2_AOI21_N3_C
x_PM_G2_AOI21_N3_Z N_Z_XI18.X0_D N_Z_XI16.X0_D N_Z_XI19.X0_D N_Z_XI17.X0_D
+ N_Z_c_170_n N_Z_c_180_n N_Z_c_174_n Z Vss PM_G2_AOI21_N3_Z
x_PM_G2_AOI21_N3_A N_A_XI18.X0_CG N_A_XI17.X0_CG N_A_c_203_n N_A_c_213_n
+ N_A_c_214_n N_A_c_204_n N_A_c_215_n N_A_c_221_n N_A_c_205_n A N_A_c_207_n Vss
+ PM_G2_AOI21_N3_A
cc_1 N_VSS_c_1_p N_VDD_c_49_n 3.30468e-19
cc_2 N_VSS_c_2_p N_VDD_c_50_n 4.89405e-19
cc_3 N_VSS_c_3_p N_VDD_c_51_n 0.00126279f
cc_4 N_VSS_c_4_p N_VDD_c_51_n 0.00161703f
cc_5 N_VSS_c_5_p N_VDD_c_51_n 2.26455e-19
cc_6 N_VSS_c_6_p N_VDD_c_51_n 0.00345242f
cc_7 N_VSS_c_7_p N_VDD_c_51_n 0.00169823f
cc_8 N_VSS_c_8_p N_VDD_c_56_n 2.74986e-19
cc_9 N_VSS_c_9_p N_VDD_c_56_n 3.26764e-19
cc_10 N_VSS_c_10_p N_VDD_c_56_n 0.00463433f
cc_11 N_VSS_c_10_p N_VDD_c_59_n 0.00166316f
cc_12 N_VSS_c_12_p N_VDD_c_60_n 4.01154e-19
cc_13 N_VSS_c_9_p N_VDD_c_61_n 0.00187494f
cc_14 N_VSS_c_14_p N_VDD_c_61_n 0.00422386f
cc_15 N_VSS_c_15_p N_VDD_c_61_n 0.00869026f
cc_16 N_VSS_c_16_p N_VDD_c_61_n 9.16632e-19
cc_17 N_VSS_c_4_p N_VDD_c_65_n 4.83895e-19
cc_18 N_VSS_c_6_p N_VDD_c_65_n 0.00105311f
cc_19 N_VSS_c_15_p N_VDD_c_65_n 0.00385589f
cc_20 N_VSS_c_15_p N_VDD_c_68_n 0.00115015f
cc_21 N_VSS_c_21_p N_B_c_105_n 3.69138e-19
cc_22 N_VSS_c_10_p N_B_c_105_n 3.72732e-19
cc_23 N_VSS_XI16.X0_PGD N_C_XI16.X0_PGS 0.00150757f
cc_24 N_VSS_c_4_p N_C_c_124_n 8.90801e-19
cc_25 N_VSS_c_5_p N_C_c_124_n 3.44698e-19
cc_26 N_VSS_c_15_p N_C_c_124_n 0.00209922f
cc_27 N_VSS_c_15_p N_C_c_127_n 5.11302e-19
cc_28 N_VSS_XI16.X0_PGD N_C_c_128_n 3.23173e-19
cc_29 N_VSS_c_3_p N_C_c_128_n 0.00480946f
cc_30 N_VSS_c_4_p N_C_c_128_n 3.44698e-19
cc_31 N_VSS_c_5_p N_C_c_128_n 6.61756e-19
cc_32 N_VSS_c_10_p N_C_c_132_n 0.00205555f
cc_33 N_VSS_c_15_p N_C_c_132_n 3.90377e-19
cc_34 N_VSS_c_34_p N_Z_c_170_n 3.43419e-19
cc_35 N_VSS_c_8_p N_Z_c_170_n 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_c_170_n 3.48267e-19
cc_37 N_VSS_c_9_p N_Z_c_170_n 3.48267e-19
cc_38 N_VSS_c_34_p N_Z_c_174_n 3.48267e-19
cc_39 N_VSS_c_8_p N_Z_c_174_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_174_n 5.71987e-19
cc_41 N_VSS_c_9_p N_Z_c_174_n 5.71987e-19
cc_42 N_VSS_c_10_p N_Z_c_174_n 3.02286e-19
cc_43 N_VSS_c_15_p N_Z_c_174_n 9.87738e-19
cc_44 N_VSS_XI16.X0_PGD N_A_c_203_n 7.5154e-19
cc_45 N_VSS_XI17.X0_PGD N_A_c_204_n 0.00163887f
cc_46 N_VSS_c_5_p N_A_c_205_n 5.05931e-19
cc_47 N_VSS_c_5_p A 2.15082e-19
cc_48 N_VSS_c_4_p N_A_c_207_n 2.15082e-19
cc_49 N_VDD_XI18.X0_PGD N_B_XI18.X0_PGS 0.00174385f
cc_50 N_VDD_c_70_p N_B_c_105_n 6.29947e-19
cc_51 N_VDD_c_71_p N_B_c_105_n 3.48267e-19
cc_52 N_VDD_XI18.X0_PGD N_B_c_110_n 3.23173e-19
cc_53 N_VDD_c_70_p N_B_c_110_n 4.44903e-19
cc_54 N_VDD_c_71_p N_B_c_110_n 6.39485e-19
cc_55 N_VDD_c_75_p N_C_XI16.X0_PGS 3.81609e-19
cc_56 N_VDD_c_76_p N_C_c_135_n 5.33384e-19
cc_57 N_VDD_c_61_n N_C_c_135_n 5.92666e-19
cc_58 N_VDD_c_51_n N_C_c_137_n 3.8746e-19
cc_59 N_VDD_XI19.X0_PGS N_C_c_138_n 8.42974e-19
cc_60 N_VDD_c_61_n N_C_c_138_n 6.25289e-19
cc_61 N_VDD_c_75_p N_C_c_124_n 0.00129723f
cc_62 N_VDD_c_50_n N_C_c_124_n 4.34459e-19
cc_63 N_VDD_c_51_n N_C_c_124_n 0.00204347f
cc_64 N_VDD_c_70_p C 2.77106e-19
cc_65 N_VDD_c_61_n C 4.49702e-19
cc_66 N_VDD_c_71_p C 2.15082e-19
cc_67 N_VDD_c_51_n N_C_c_127_n 5.0979e-19
cc_68 N_VDD_c_75_p N_C_c_128_n 3.66936e-19
cc_69 N_VDD_c_51_n N_C_c_128_n 2.64932e-19
cc_70 N_VDD_c_90_p N_Z_c_180_n 3.43419e-19
cc_71 N_VDD_c_91_p N_Z_c_180_n 3.43419e-19
cc_72 N_VDD_c_50_n N_Z_c_180_n 3.72199e-19
cc_73 N_VDD_c_51_n N_Z_c_180_n 2.74986e-19
cc_74 N_VDD_c_60_n N_Z_c_180_n 3.72199e-19
cc_75 N_VDD_c_90_p N_Z_c_174_n 3.48267e-19
cc_76 N_VDD_c_91_p N_Z_c_174_n 3.48267e-19
cc_77 N_VDD_c_50_n N_Z_c_174_n 5.09542e-19
cc_78 N_VDD_c_51_n N_Z_c_174_n 5.72568e-19
cc_79 N_VDD_c_60_n N_Z_c_174_n 7.72285e-19
cc_80 N_VDD_c_61_n N_Z_c_174_n 0.00179861f
cc_81 N_VDD_XI18.X0_PGD N_A_c_203_n 6.25166e-19
cc_82 N_VDD_XI19.X0_PGD N_A_c_204_n 3.70201e-19
cc_83 N_VDD_c_61_n A 4.8807e-19
cc_84 N_VDD_c_61_n N_A_c_207_n 3.66936e-19
cc_85 N_B_c_113_p N_C_XI16.X0_PGS 0.0020206f
cc_86 N_B_XI18.X0_PGS N_C_XI19.X0_CG 2.46172e-19
cc_87 N_B_c_113_p N_C_XI17.X0_PGS 4.66827e-19
cc_88 N_B_c_105_n N_C_c_132_n 2.19701e-19
cc_89 N_B_XI18.X0_PGS N_Z_c_174_n 2.61881e-19
cc_90 N_B_XI18.X0_PGS N_A_XI18.X0_CG 0.00881601f
cc_91 N_B_c_113_p N_A_c_213_n 0.00191565f
cc_92 N_B_XI18.X0_PGS N_A_c_214_n 6.07734e-19
cc_93 N_B_c_113_p N_A_c_215_n 0.00136534f
cc_94 N_B_c_113_p N_A_c_207_n 2.87722e-19
cc_95 N_C_c_135_n N_Z_c_174_n 9.83688e-19
cc_96 N_C_c_124_n N_Z_c_174_n 0.00308891f
cc_97 C N_Z_c_174_n 0.00140888f
cc_98 N_C_c_127_n N_Z_c_174_n 0.00195497f
cc_99 N_C_c_132_n N_Z_c_174_n 2.70867e-19
cc_100 N_C_XI19.X0_CG N_A_XI18.X0_CG 5.48933e-19
cc_101 N_C_c_135_n N_A_XI18.X0_CG 5.60239e-19
cc_102 N_C_XI17.X0_PGS N_A_c_203_n 8.10159e-19
cc_103 N_C_c_138_n N_A_c_203_n 0.00121323f
cc_104 N_C_XI17.X0_PGS N_A_c_221_n 4.42555e-19
cc_105 N_C_c_135_n N_A_c_205_n 9.47282e-19
cc_106 N_C_c_135_n A 4.56568e-19
cc_107 C A 6.3743e-19
cc_108 N_C_XI17.X0_PGS N_A_c_207_n 0.00570455f
cc_109 N_C_c_135_n N_A_c_207_n 6.1245e-19
cc_110 N_C_c_138_n N_A_c_207_n 0.00239404f
cc_111 C N_A_c_207_n 4.56568e-19
cc_112 N_Z_c_174_n N_A_XI18.X0_CG 5.52516e-19
cc_113 N_Z_c_170_n N_A_c_203_n 3.56294e-19
cc_114 N_Z_c_174_n N_A_c_203_n 3.092e-19
cc_115 N_Z_c_180_n N_A_c_215_n 5.66216e-19
cc_116 N_Z_c_174_n A 0.00149422f
cc_117 N_Z_c_174_n N_A_c_207_n 9.53426e-19
*
.ends
*
*
.subckt AOI21_HPNW12 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 B0 Y A0) G2_AOI21_N3
.ends
*
* File: G2_BUF1_N3.pex.netlist
* Created: Wed Mar  2 15:50:41 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_BUF1_N3_VDD 2 4 7 11 28 30 32 44 48 52 54 56 57 61 65 67 71 75 78
+ 90 95 Vss
c55 95 Vss 0.00494983f
c56 90 Vss 0.00475556f
c57 80 Vss 9.22237e-19
c58 79 Vss 9.22237e-19
c59 75 Vss 0.00138508f
c60 71 Vss 9.81533e-19
c61 68 Vss 0.00177515f
c62 67 Vss 0.00751016f
c63 65 Vss 0.0012592f
c64 61 Vss 0.0012592f
c65 57 Vss 0.00744668f
c66 56 Vss 0.00466777f
c67 54 Vss 0.00779694f
c68 52 Vss 0.00466777f
c69 51 Vss 0.00177515f
c70 48 Vss 0.00810125f
c71 44 Vss 0.0100206f
c72 32 Vss 0.0356247f
c73 31 Vss 0.102427f
c74 28 Vss 0.0356247f
c75 27 Vss 0.102427f
c76 11 Vss 0.378484f
c77 7 Vss 0.378484f
r78 75 95 1.16709
r79 73 75 2.16729
r80 71 90 1.16709
r81 69 71 2.16729
r82 67 73 0.652036
r83 67 68 10.1279
r84 63 80 0.0828784
r85 63 65 1.82344
r86 59 79 0.0828784
r87 59 61 1.82344
r88 58 78 0.326018
r89 57 69 0.652036
r90 57 58 10.1279
r91 56 68 0.652036
r92 55 80 0.551426
r93 55 56 5.50157
r94 54 80 0.551426
r95 53 79 0.551426
r96 53 54 8.58579
r97 52 79 0.551426
r98 51 78 0.326018
r99 51 52 5.50157
r100 48 65 1.16709
r101 44 61 1.16709
r102 34 95 0.0476429
r103 32 34 1.45875
r104 31 38 0.652036
r105 31 34 1.45875
r106 30 90 0.0476429
r107 28 30 1.45875
r108 27 35 0.652036
r109 27 30 1.45875
r110 24 32 0.652036
r111 21 28 0.652036
r112 11 38 5.1348
r113 11 24 5.1348
r114 7 35 5.1348
r115 7 21 5.1348
r116 4 48 0.123773
r117 2 44 0.123773
.ends

.subckt PM_G2_BUF1_N3_VSS 3 7 10 12 27 28 31 32 45 49 52 57 62 67 72 77 97 98 99
+ 100 101 105 110 112 114 116 Vss
c52 118 Vss 6.78504e-19
c53 117 Vss 6.78504e-19
c54 114 Vss 0.00360796f
c55 112 Vss 0.00582053f
c56 110 Vss 0.00360796f
c57 109 Vss 0.0013648f
c58 105 Vss 0.0010737f
c59 101 Vss 9.14356e-19
c60 100 Vss 5.83649e-19
c61 99 Vss 0.00682958f
c62 98 Vss 5.83649e-19
c63 97 Vss 0.00550031f
c64 77 Vss 0.00392669f
c65 72 Vss 0.00392498f
c66 67 Vss 1.62518e-19
c67 62 Vss 7.10513e-22
c68 57 Vss 8.49747e-19
c69 52 Vss 0.00100529f
c70 49 Vss 0.0100686f
c71 45 Vss 0.00814922f
c72 32 Vss 0.0350852f
c73 31 Vss 0.0994129f
c74 28 Vss 0.0350852f
c75 27 Vss 0.0994129f
c76 7 Vss 0.377694f
c77 3 Vss 0.377694f
r78 113 118 0.551426
r79 113 114 5.50157
r80 112 118 0.551426
r81 111 117 0.551426
r82 111 112 8.58579
r83 110 117 0.551426
r84 109 116 0.326018
r85 109 110 5.50157
r86 105 118 0.0828784
r87 101 117 0.0828784
r88 99 114 0.652036
r89 99 100 10.1279
r90 97 116 0.326018
r91 97 98 10.1279
r92 93 100 0.652036
r93 89 98 0.652036
r94 67 105 1.82344
r95 62 101 1.82344
r96 57 77 1.16709
r97 57 93 2.16729
r98 52 72 1.16709
r99 52 89 2.16729
r100 49 67 1.16709
r101 45 62 1.16709
r102 34 77 0.0476429
r103 32 34 1.45875
r104 31 38 0.652036
r105 31 34 1.45875
r106 30 72 0.0476429
r107 28 30 1.45875
r108 27 35 0.652036
r109 27 30 1.45875
r110 24 32 0.652036
r111 21 28 0.652036
r112 12 49 0.123773
r113 10 45 0.123773
r114 7 38 5.1348
r115 7 24 5.1348
r116 3 35 5.1348
r117 3 21 5.1348
.ends

.subckt PM_G2_BUF1_N3_A 2 4 12 24 27 Vss
c13 27 Vss 0.00315166f
c14 24 Vss 1.56823e-19
c15 12 Vss 0.20431f
c16 9 Vss 0.180512f
c17 7 Vss 0.0247918f
c18 4 Vss 0.193588f
r19 24 27 1.16709
r20 15 27 0.0476429
r21 13 15 0.326018
r22 13 15 0.1167
r23 12 16 0.652036
r24 12 15 6.7686
r25 9 27 0.357321
r26 7 15 0.326018
r27 7 9 0.40845
r28 4 16 5.1348
r29 2 9 4.72635
.ends

.subckt PM_G2_BUF1_N3_Z 2 4 13 16 19 Vss
c13 16 Vss 3.73795e-19
c14 13 Vss 0.00513911f
c15 4 Vss 0.00176592f
r16 16 19 0.0416786
r17 13 16 1.16709
r18 4 13 0.123773
r19 2 13 0.123773
.ends

.subckt PM_G2_BUF1_N3_NET17 2 4 6 8 18 33 36 41 50 58 Vss
c31 58 Vss 5.10694e-19
c32 50 Vss 0.0034988f
c33 41 Vss 0.0021514f
c34 36 Vss 0.0018043f
c35 33 Vss 0.00513911f
c36 22 Vss 0.0247918f
c37 19 Vss 0.0299669f
c38 18 Vss 0.173331f
c39 8 Vss 0.00176592f
c40 6 Vss 0.180667f
c41 2 Vss 0.192541f
r42 54 58 0.653045
r43 41 50 1.16709
r44 41 58 2.1395
r45 36 54 5.29318
r46 33 36 1.16709
r47 28 50 0.0476429
r48 26 50 0.357321
r49 22 28 0.326018
r50 22 26 0.40845
r51 19 28 6.7686
r52 18 28 0.326018
r53 18 28 0.1167
r54 15 19 0.652036
r55 8 33 0.123773
r56 6 26 4.72635
r57 4 33 0.123773
r58 2 15 5.1348
.ends

.subckt G2_BUF1_N3  VDD VSS A Z
*
* Z	Z
* A	A
* VSS	VSS
* VDD	VDD
XI14.X0 N_Z_XI14.X0_D N_VSS_XI14.X0_PGD N_NET17_XI14.X0_CG N_VSS_XI14.X0_PGD
+ N_VDD_XI14.X0_S TIGFET_HPNW12
XI11.X0 N_NET17_XI11.X0_D N_VSS_XI11.X0_PGD N_A_XI11.X0_CG N_VSS_XI11.X0_PGD
+ N_VDD_XI11.X0_S TIGFET_HPNW12
XI13.X0 N_Z_XI13.X0_D N_VDD_XI13.X0_PGD N_NET17_XI13.X0_CG N_VDD_XI13.X0_PGD
+ N_VSS_XI13.X0_S TIGFET_HPNW12
XI12.X0 N_NET17_XI12.X0_D N_VDD_XI12.X0_PGD N_A_XI12.X0_CG N_VDD_XI12.X0_PGD
+ N_VSS_XI12.X0_S TIGFET_HPNW12
*
x_PM_G2_BUF1_N3_VDD N_VDD_XI14.X0_S N_VDD_XI11.X0_S N_VDD_XI13.X0_PGD
+ N_VDD_XI12.X0_PGD N_VDD_c_4_p N_VDD_c_50_p N_VDD_c_8_p N_VDD_c_36_p
+ N_VDD_c_45_p N_VDD_c_6_p N_VDD_c_34_p N_VDD_c_3_p N_VDD_c_5_p N_VDD_c_38_p
+ N_VDD_c_46_p N_VDD_c_9_p N_VDD_c_13_p N_VDD_c_17_p VDD N_VDD_c_14_p
+ N_VDD_c_18_p Vss PM_G2_BUF1_N3_VDD
x_PM_G2_BUF1_N3_VSS N_VSS_XI14.X0_PGD N_VSS_XI11.X0_PGD N_VSS_XI13.X0_S
+ N_VSS_XI12.X0_S N_VSS_c_59_n N_VSS_c_61_n N_VSS_c_63_n N_VSS_c_65_n
+ N_VSS_c_93_p N_VSS_c_99_p N_VSS_c_66_n N_VSS_c_70_n N_VSS_c_94_p N_VSS_c_100_p
+ N_VSS_c_74_n N_VSS_c_78_n N_VSS_c_81_n N_VSS_c_82_n N_VSS_c_83_n N_VSS_c_84_n
+ N_VSS_c_96_p N_VSS_c_103_p N_VSS_c_85_n N_VSS_c_104_p N_VSS_c_86_n VSS Vss
+ PM_G2_BUF1_N3_VSS
x_PM_G2_BUF1_N3_A N_A_XI11.X0_CG N_A_XI12.X0_CG N_A_c_108_n A N_A_c_111_n Vss
+ PM_G2_BUF1_N3_A
x_PM_G2_BUF1_N3_Z N_Z_XI14.X0_D N_Z_XI13.X0_D N_Z_c_121_n N_Z_c_124_n Z Vss
+ PM_G2_BUF1_N3_Z
x_PM_G2_BUF1_N3_NET17 N_NET17_XI14.X0_CG N_NET17_XI11.X0_D N_NET17_XI13.X0_CG
+ N_NET17_XI12.X0_D N_NET17_c_135_n N_NET17_c_137_n N_NET17_c_139_n
+ N_NET17_c_142_n N_NET17_c_146_n N_NET17_c_147_n Vss PM_G2_BUF1_N3_NET17
cc_1 N_VDD_XI13.X0_PGD N_VSS_XI14.X0_PGD 0.00200662f
cc_2 N_VDD_XI12.X0_PGD N_VSS_XI11.X0_PGD 0.00200662f
cc_3 N_VDD_c_3_p N_VSS_XI11.X0_PGD 4.00543e-19
cc_4 N_VDD_c_4_p N_VSS_c_59_n 0.00200662f
cc_5 N_VDD_c_5_p N_VSS_c_59_n 3.89167e-19
cc_6 N_VDD_c_6_p N_VSS_c_61_n 4.00543e-19
cc_7 N_VDD_c_5_p N_VSS_c_61_n 4.0633e-19
cc_8 N_VDD_c_8_p N_VSS_c_63_n 0.00200662f
cc_9 N_VDD_c_9_p N_VSS_c_63_n 3.89167e-19
cc_10 N_VDD_c_9_p N_VSS_c_65_n 4.0633e-19
cc_11 N_VDD_c_6_p N_VSS_c_66_n 9.94764e-19
cc_12 N_VDD_c_5_p N_VSS_c_66_n 0.00162079f
cc_13 N_VDD_c_13_p N_VSS_c_66_n 0.00106273f
cc_14 N_VDD_c_14_p N_VSS_c_66_n 3.48267e-19
cc_15 N_VDD_c_3_p N_VSS_c_70_n 9.94764e-19
cc_16 N_VDD_c_9_p N_VSS_c_70_n 0.00141604f
cc_17 N_VDD_c_17_p N_VSS_c_70_n 0.00110056f
cc_18 N_VDD_c_18_p N_VSS_c_70_n 3.48267e-19
cc_19 N_VDD_c_6_p N_VSS_c_74_n 3.66936e-19
cc_20 N_VDD_c_5_p N_VSS_c_74_n 2.2543e-19
cc_21 N_VDD_c_13_p N_VSS_c_74_n 3.99794e-19
cc_22 N_VDD_c_14_p N_VSS_c_74_n 6.489e-19
cc_23 N_VDD_c_3_p N_VSS_c_78_n 3.66936e-19
cc_24 N_VDD_c_9_p N_VSS_c_78_n 0.00114409f
cc_25 N_VDD_c_18_p N_VSS_c_78_n 6.489e-19
cc_26 N_VDD_c_5_p N_VSS_c_81_n 0.00589548f
cc_27 N_VDD_c_5_p N_VSS_c_82_n 0.0017359f
cc_28 N_VDD_c_9_p N_VSS_c_83_n 0.00593021f
cc_29 N_VDD_c_9_p N_VSS_c_84_n 0.0017359f
cc_30 N_VDD_c_13_p N_VSS_c_85_n 3.85245e-19
cc_31 N_VDD_c_17_p N_VSS_c_86_n 3.85245e-19
cc_32 N_VDD_XI13.X0_PGD N_A_c_108_n 4.14544e-19
cc_33 N_VDD_XI12.X0_PGD N_A_c_108_n 4.09718e-19
cc_34 N_VDD_c_34_p A 9.3432e-19
cc_35 N_VDD_c_34_p N_A_c_111_n 5.79991e-19
cc_36 N_VDD_c_36_p N_Z_c_121_n 3.43419e-19
cc_37 N_VDD_c_5_p N_Z_c_121_n 2.74986e-19
cc_38 N_VDD_c_38_p N_Z_c_121_n 3.72199e-19
cc_39 N_VDD_c_36_p N_Z_c_124_n 3.48267e-19
cc_40 N_VDD_c_5_p N_Z_c_124_n 3.66281e-19
cc_41 N_VDD_c_38_p N_Z_c_124_n 7.4527e-19
cc_42 N_VDD_c_34_p N_NET17_XI14.X0_CG 3.93898e-19
cc_43 N_VDD_XI13.X0_PGD N_NET17_c_135_n 4.09718e-19
cc_44 N_VDD_XI12.X0_PGD N_NET17_c_135_n 4.14544e-19
cc_45 N_VDD_c_45_p N_NET17_c_137_n 3.43419e-19
cc_46 N_VDD_c_46_p N_NET17_c_137_n 3.72199e-19
cc_47 N_VDD_c_45_p N_NET17_c_139_n 3.48267e-19
cc_48 N_VDD_c_46_p N_NET17_c_139_n 8.0086e-19
cc_49 N_VDD_c_9_p N_NET17_c_139_n 3.21336e-19
cc_50 N_VDD_c_50_p N_NET17_c_142_n 2.21762e-19
cc_51 N_VDD_c_34_p N_NET17_c_142_n 2.74452e-19
cc_52 N_VDD_c_13_p N_NET17_c_142_n 2.88301e-19
cc_53 N_VDD_c_14_p N_NET17_c_142_n 2.30774e-19
cc_54 N_VDD_c_13_p N_NET17_c_146_n 2.28697e-19
cc_55 N_VDD_c_34_p N_NET17_c_147_n 7.45369e-19
cc_56 N_VSS_XI14.X0_PGD N_A_c_108_n 4.14544e-19
cc_57 N_VSS_XI11.X0_PGD N_A_c_108_n 4.09718e-19
cc_58 N_VSS_c_66_n A 2.26871e-19
cc_59 N_VSS_c_70_n A 3.35067e-19
cc_60 N_VSS_c_78_n A 2.30774e-19
cc_61 N_VSS_c_70_n N_A_c_111_n 2.28892e-19
cc_62 N_VSS_c_93_p N_Z_c_121_n 3.43419e-19
cc_63 N_VSS_c_94_p N_Z_c_121_n 3.48267e-19
cc_64 N_VSS_c_94_p N_Z_c_124_n 5.37696e-19
cc_65 N_VSS_c_96_p N_Z_c_124_n 2.7826e-19
cc_66 N_VSS_XI14.X0_PGD N_NET17_c_135_n 4.09718e-19
cc_67 N_VSS_XI11.X0_PGD N_NET17_c_135_n 4.14544e-19
cc_68 N_VSS_c_99_p N_NET17_c_137_n 3.43419e-19
cc_69 N_VSS_c_100_p N_NET17_c_137_n 3.48267e-19
cc_70 N_VSS_c_100_p N_NET17_c_139_n 4.8288e-19
cc_71 N_VSS_c_83_n N_NET17_c_139_n 3.94979e-19
cc_72 N_VSS_c_103_p N_NET17_c_139_n 5.49885e-19
cc_73 N_VSS_c_104_p N_NET17_c_139_n 0.00142716f
cc_74 N_VSS_c_104_p N_NET17_c_142_n 0.00119345f
cc_75 N_VSS_c_81_n N_NET17_c_147_n 6.75516e-19
cc_76 N_VSS_c_83_n N_NET17_c_147_n 4.01006e-19
cc_77 N_A_c_108_n N_NET17_c_135_n 0.00945061f
cc_78 N_A_c_108_n N_NET17_c_137_n 4.98287e-19
cc_79 A N_NET17_c_139_n 8.54729e-19
cc_80 N_Z_c_121_n N_NET17_c_135_n 4.98287e-19
cc_81 N_Z_c_121_n N_NET17_c_137_n 3.80999e-19
cc_82 N_Z_c_124_n N_NET17_c_147_n 2.07279e-19
*
.ends
*
*
.subckt BUF1_HPNW12 A Y VDD VSS
xgate (VDD VSS A Y) G2_BUF1_N3
.ends
*
* File: G3_DFFQ1_N3.pex.netlist
* Created: Wed Apr  6 11:25:19 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_DFFQ1_N3_VSS 2 4 6 8 10 12 14 29 42 44 49 55 59 64 67 72 78 83 88
+ 93 102 111 117 126 127 128 129 133 138 143 149 155 157 162 164 166 167 168 Vss
c101 168 Vss 4.28045e-19
c102 167 Vss 3.75522e-19
c103 166 Vss 3.75522e-19
c104 165 Vss 6.20041e-19
c105 164 Vss 0.00614697f
c106 162 Vss 0.00220014f
c107 157 Vss 0.0014078f
c108 155 Vss 0.00256807f
c109 149 Vss 0.00450029f
c110 143 Vss 0.00309494f
c111 133 Vss 0.00200475f
c112 129 Vss 6.50617e-19
c113 128 Vss 8.16747e-19
c114 127 Vss 0.00572724f
c115 126 Vss 0.0020774f
c116 117 Vss 0.00492488f
c117 111 Vss 0.00403629f
c118 102 Vss 0.00419844f
c119 93 Vss 2.01624e-19
c120 88 Vss 9.8978e-19
c121 83 Vss 8.45647e-19
c122 78 Vss 0.00151704f
c123 72 Vss 0.0130885f
c124 67 Vss 0.00136241f
c125 64 Vss 0.0111802f
c126 59 Vss 0.00964026f
c127 55 Vss 0.00801889f
c128 49 Vss 0.0568987f
c129 44 Vss 0.0568992f
c130 42 Vss 8.92801e-20
c131 29 Vss 0.0356247f
c132 28 Vss 0.101312f
c133 14 Vss 0.189842f
c134 8 Vss 0.191315f
c135 6 Vss 0.188337f
c136 4 Vss 0.188444f
r137 163 168 0.551426
r138 163 164 18.3386
r139 162 168 0.551426
r140 161 162 5.54325
r141 157 168 0.0828784
r142 156 167 0.494161
r143 155 164 0.652036
r144 155 156 4.37625
r145 151 167 0.128424
r146 150 166 0.494161
r147 149 161 0.652036
r148 149 150 10.1279
r149 145 166 0.128424
r150 144 165 0.494161
r151 143 167 0.494161
r152 143 144 7.46046
r153 139 165 0.128424
r154 133 165 0.494161
r155 133 138 1.00029
r156 127 166 0.494161
r157 127 128 15.8795
r158 126 129 0.655813
r159 125 128 0.652036
r160 125 126 5.54325
r161 111 114 0.05
r162 93 157 1.82344
r163 88 117 1.16709
r164 88 151 2.16729
r165 83 114 1.16709
r166 83 145 2.20896
r167 78 139 6.16843
r168 75 138 1.29204
r169 72 102 1.16709
r170 72 75 15.5878
r171 67 129 1.82344
r172 64 93 1.16709
r173 59 78 1.16709
r174 55 67 1.16709
r175 49 117 0.197068
r176 46 49 1.2837
r177 42 111 0.197068
r178 42 44 1.2837
r179 38 46 0.0685365
r180 35 44 0.0685365
r181 31 102 0.0476429
r182 29 31 1.45875
r183 28 32 0.652036
r184 28 31 1.45875
r185 25 29 0.652036
r186 14 38 5.1348
r187 12 64 0.123773
r188 10 59 0.123773
r189 8 35 5.1348
r190 6 32 5.1348
r191 4 25 5.1348
r192 2 55 0.123773
.ends

.subckt PM_G3_DFFQ1_N3_CK 2 4 6 8 18 21 25 35 41 Vss
c33 41 Vss 0.00492267f
c34 35 Vss 3.25681e-19
c35 33 Vss 0.0299314f
c36 25 Vss 0.166167f
c37 21 Vss 8.92801e-20
c38 18 Vss 0.18663f
c39 15 Vss 0.180502f
c40 13 Vss 0.0247918f
c41 6 Vss 0.659388f
c42 4 Vss 0.191169f
r43 41 44 0.05
r44 38 44 1.16709
r45 35 38 0.0416786
r46 26 33 0.494161
r47 25 27 0.652036
r48 25 26 4.84305
r49 22 33 0.128424
r50 21 41 0.0238214
r51 19 21 0.326018
r52 19 21 0.1167
r53 18 33 0.494161
r54 18 21 6.7686
r55 15 41 0.357321
r56 13 21 0.326018
r57 13 15 0.3501
r58 6 8 17.9718
r59 6 27 5.1348
r60 4 22 5.1348
r61 2 15 4.7847
.ends

.subckt PM_G3_DFFQ1_N3_VDD 2 4 6 8 10 12 14 28 42 44 49 56 60 63 64 65 70 72 76
+ 78 79 82 84 86 91 93 95 96 98 99 100 102 104 113 118 Vss
c107 118 Vss 0.00533757f
c108 113 Vss 0.00573314f
c109 104 Vss 0.00489453f
c110 100 Vss 4.52364e-19
c111 99 Vss 2.39889e-19
c112 98 Vss 4.43992e-19
c113 96 Vss 0.00375805f
c114 95 Vss 4.90076e-19
c115 93 Vss 0.00385631f
c116 91 Vss 0.0108071f
c117 86 Vss 0.00177107f
c118 84 Vss 0.0031515f
c119 82 Vss 0.00100814f
c120 79 Vss 4.90412e-19
c121 78 Vss 0.00546064f
c122 76 Vss 6.46297e-19
c123 72 Vss 0.00354521f
c124 70 Vss 0.00226527f
c125 67 Vss 0.00183337f
c126 65 Vss 8.65196e-19
c127 64 Vss 0.00754197f
c128 63 Vss 0.00697044f
c129 60 Vss 0.0112146f
c130 56 Vss 0.0070753f
c131 49 Vss 0.0589116f
c132 44 Vss 0.0581535f
c133 42 Vss 7.85965e-20
c134 29 Vss 0.0372509f
c135 28 Vss 0.101007f
c136 12 Vss 0.191734f
c137 10 Vss 0.189852f
c138 8 Vss 0.00143493f
c139 4 Vss 0.190684f
c140 2 Vss 0.189513f
r141 118 121 0.05
r142 95 104 1.16709
r143 95 96 0.470345
r144 93 102 0.326018
r145 92 100 0.551426
r146 92 93 5.50157
r147 91 100 0.551426
r148 90 91 18.3803
r149 86 100 0.0828784
r150 86 88 1.82344
r151 85 99 0.494161
r152 84 90 0.652036
r153 84 85 4.37625
r154 82 121 1.16709
r155 80 99 0.128424
r156 80 82 2.20896
r157 78 102 0.326018
r158 78 79 10.1279
r159 76 113 1.16709
r160 74 79 0.652036
r161 74 76 2.16729
r162 73 98 0.494161
r163 72 99 0.494161
r164 72 73 7.46046
r165 68 98 0.128424
r166 68 70 6.21011
r167 67 96 3.82922
r168 64 98 0.494161
r169 64 65 13.0037
r170 63 67 0.655813
r171 62 65 0.652036
r172 62 63 10.2113
r173 60 88 1.16709
r174 56 70 1.16709
r175 49 118 0.197068
r176 46 49 1.2837
r177 42 113 0.197068
r178 42 44 1.2837
r179 38 46 0.0685365
r180 35 44 0.0685365
r181 31 104 0.0476429
r182 29 31 1.45875
r183 28 32 0.652036
r184 28 31 1.45875
r185 25 29 0.652036
r186 14 60 0.123773
r187 12 38 5.1348
r188 10 35 5.1348
r189 8 56 0.123773
r190 6 56 0.123773
r191 4 25 5.1348
r192 2 32 5.1348
.ends

.subckt PM_G3_DFFQ1_N3_CKN 2 4 6 8 18 25 28 33 50 Vss
c37 51 Vss 0.00128789f
c38 50 Vss 0.00701318f
c39 33 Vss 3.33899e-19
c40 28 Vss 0.00179767f
c41 25 Vss 0.00520172f
c42 18 Vss 7.22113e-19
c43 6 Vss 0.584002f
c44 4 Vss 0.00143493f
r45 50 51 14.6709
r46 46 51 0.652036
r47 33 50 0.531835
r48 28 46 5.835
r49 25 28 1.16709
r50 18 33 1.16709
r51 8 18 8.9859
r52 6 18 8.9859
r53 4 25 0.123773
r54 2 25 0.123773
.ends

.subckt PM_G3_DFFQ1_N3_D 2 4 11 12 22 25 28 Vss
c24 28 Vss 0.00196994f
c25 25 Vss 4.67436e-19
c26 12 Vss 0.214507f
c27 11 Vss 8.44702e-20
c28 7 Vss 0.0247918f
c29 4 Vss 0.191884f
c30 2 Vss 0.180391f
r31 25 28 1.16709
r32 22 25 0.0364688
r33 15 28 0.0476429
r34 13 15 0.326018
r35 13 15 0.1167
r36 12 16 0.652036
r37 12 15 6.7686
r38 11 28 0.357321
r39 7 15 0.326018
r40 7 11 0.40845
r41 4 16 5.1348
r42 2 11 4.72635
.ends

.subckt PM_G3_DFFQ1_N3_X 2 4 6 8 17 20 23 33 35 39 41 47 Vss
c46 47 Vss 0.00165819f
c47 41 Vss 5.1586e-19
c48 39 Vss 0.00126373f
c49 35 Vss 0.00198822f
c50 33 Vss 0.00525025f
c51 23 Vss 7.81442e-20
c52 20 Vss 0.214848f
c53 17 Vss 0.180344f
c54 15 Vss 0.0247918f
c55 8 Vss 0.191809f
c56 6 Vss 0.00143493f
r57 44 47 1.16709
r58 41 44 2.08393
r59 37 39 6.16843
r60 36 41 0.0685365
r61 35 37 0.652036
r62 35 36 1.70882
r63 33 39 1.16709
r64 23 47 0.0476429
r65 21 23 0.326018
r66 21 23 0.1167
r67 20 24 0.652036
r68 20 23 6.7686
r69 17 47 0.357321
r70 15 23 0.326018
r71 15 17 0.40845
r72 8 24 5.1348
r73 6 33 0.123773
r74 4 17 4.72635
r75 2 33 0.123773
.ends

.subckt PM_G3_DFFQ1_N3_Q 2 4 13 16 Vss
c12 16 Vss 3.46649e-19
c13 13 Vss 0.0045421f
c14 4 Vss 0.00143493f
r15 16 19 0.0416786
r16 13 19 1.16709
r17 4 13 0.123773
r18 2 13 0.123773
.ends

.subckt G3_DFFQ1_N3  VSS CK VDD D Q
*
* Q	Q
* D	D
* VDD	VDD
* CK	CK
* VSS	VSS
XI0.X0 N_CKN_XI0.X0_D N_VDD_XI0.X0_PGD N_CK_XI0.X0_CG N_VDD_XI0.X0_PGS
+ N_VSS_XI0.X0_S TIGFET_HPNW12
XI1.X0 N_CKN_XI1.X0_D N_VSS_XI1.X0_PGD N_CK_XI1.X0_CG N_VSS_XI1.X0_PGS
+ N_VDD_XI1.X0_S TIGFET_HPNW12
XI13.X0 N_X_XI13.X0_D N_VSS_XI13.X0_PGD N_D_XI13.X0_CG N_CK_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW12
XI4.X0 N_Q_XI4.X0_D N_VDD_XI4.X0_PGD N_X_XI4.X0_CG N_CK_XI4.X0_PGS
+ N_VSS_XI4.X0_S TIGFET_HPNW12
XI12.X0 N_X_XI12.X0_D N_VDD_XI12.X0_PGD N_D_XI12.X0_CG N_CKN_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW12
XI5.X0 N_Q_XI5.X0_D N_VSS_XI5.X0_PGD N_X_XI5.X0_CG N_CKN_XI5.X0_PGS
+ N_VDD_XI5.X0_S TIGFET_HPNW12
*
x_PM_G3_DFFQ1_N3_VSS N_VSS_XI0.X0_S N_VSS_XI1.X0_PGD N_VSS_XI1.X0_PGS
+ N_VSS_XI13.X0_PGD N_VSS_XI4.X0_S N_VSS_XI12.X0_S N_VSS_XI5.X0_PGD N_VSS_c_11_p
+ N_VSS_c_81_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_14_p N_VSS_c_99_p N_VSS_c_41_p
+ N_VSS_c_15_p N_VSS_c_3_p N_VSS_c_30_p N_VSS_c_21_p N_VSS_c_31_p N_VSS_c_42_p
+ N_VSS_c_54_p N_VSS_c_4_p N_VSS_c_34_p N_VSS_c_16_p N_VSS_c_7_p N_VSS_c_20_p
+ N_VSS_c_17_p N_VSS_c_78_p VSS N_VSS_c_35_p N_VSS_c_27_p N_VSS_c_36_p
+ N_VSS_c_44_p N_VSS_c_46_p N_VSS_c_47_p N_VSS_c_28_p N_VSS_c_37_p N_VSS_c_48_p
+ Vss PM_G3_DFFQ1_N3_VSS
x_PM_G3_DFFQ1_N3_CK N_CK_XI0.X0_CG N_CK_XI1.X0_CG N_CK_XI13.X0_PGS
+ N_CK_XI4.X0_PGS N_CK_c_106_n N_CK_c_124_p N_CK_c_107_n CK N_CK_c_114_p Vss
+ PM_G3_DFFQ1_N3_CK
x_PM_G3_DFFQ1_N3_VDD N_VDD_XI0.X0_PGD N_VDD_XI0.X0_PGS N_VDD_XI1.X0_S
+ N_VDD_XI13.X0_S N_VDD_XI4.X0_PGD N_VDD_XI12.X0_PGD N_VDD_XI5.X0_S
+ N_VDD_c_138_n N_VDD_c_224_p N_VDD_c_139_n N_VDD_c_140_n N_VDD_c_197_n
+ N_VDD_c_236_p N_VDD_c_141_n N_VDD_c_145_n N_VDD_c_147_n N_VDD_c_148_n
+ N_VDD_c_150_n N_VDD_c_156_n N_VDD_c_159_n N_VDD_c_165_n N_VDD_c_166_n
+ N_VDD_c_168_n N_VDD_c_171_n N_VDD_c_172_n N_VDD_c_176_n N_VDD_c_180_n
+ N_VDD_c_182_n N_VDD_c_184_n N_VDD_c_185_n N_VDD_c_186_n VDD N_VDD_c_187_n
+ N_VDD_c_189_n N_VDD_c_192_n Vss PM_G3_DFFQ1_N3_VDD
x_PM_G3_DFFQ1_N3_CKN N_CKN_XI0.X0_D N_CKN_XI1.X0_D N_CKN_XI12.X0_PGS
+ N_CKN_XI5.X0_PGS N_CKN_c_257_n N_CKN_c_242_n N_CKN_c_244_n N_CKN_c_248_n
+ N_CKN_c_249_n Vss PM_G3_DFFQ1_N3_CKN
x_PM_G3_DFFQ1_N3_D N_D_XI13.X0_CG N_D_XI12.X0_CG N_D_c_279_n N_D_c_280_n D
+ N_D_c_281_n N_D_c_284_n Vss PM_G3_DFFQ1_N3_D
x_PM_G3_DFFQ1_N3_X N_X_XI13.X0_D N_X_XI4.X0_CG N_X_XI12.X0_D N_X_XI5.X0_CG
+ N_X_c_314_n N_X_c_303_n N_X_c_317_n N_X_c_304_n N_X_c_330_n N_X_c_306_n
+ N_X_c_310_n N_X_c_312_n Vss PM_G3_DFFQ1_N3_X
x_PM_G3_DFFQ1_N3_Q N_Q_XI4.X0_D N_Q_XI5.X0_D N_Q_c_349_n Q Vss PM_G3_DFFQ1_N3_Q
cc_1 N_VSS_XI1.X0_PGS N_CK_XI13.X0_PGS 0.00316278f
cc_2 N_VSS_XI13.X0_PGD N_CK_XI13.X0_PGS 0.00164185f
cc_3 N_VSS_c_3_p N_CK_XI13.X0_PGS 8.34822e-19
cc_4 N_VSS_c_4_p N_CK_XI13.X0_PGS 4.02129e-19
cc_5 N_VSS_XI1.X0_PGD N_CK_c_106_n 4.20343e-19
cc_6 N_VSS_XI1.X0_PGS N_CK_c_107_n 4.31283e-19
cc_7 N_VSS_c_7_p CK 5.33707e-19
cc_8 N_VSS_XI1.X0_PGD N_VDD_XI0.X0_PGD 0.00196344f
cc_9 N_VSS_XI5.X0_PGD N_VDD_XI4.X0_PGD 0.00221489f
cc_10 N_VSS_XI13.X0_PGD N_VDD_XI12.X0_PGD 0.00211593f
cc_11 N_VSS_c_11_p N_VDD_c_138_n 0.00196344f
cc_12 N_VSS_c_12_p N_VDD_c_139_n 0.00221489f
cc_13 N_VSS_c_13_p N_VDD_c_140_n 0.00211593f
cc_14 N_VSS_c_14_p N_VDD_c_141_n 9.5668e-19
cc_15 N_VSS_c_15_p N_VDD_c_141_n 0.00165395f
cc_16 N_VSS_c_16_p N_VDD_c_141_n 0.00423852f
cc_17 N_VSS_c_17_p N_VDD_c_141_n 0.00186049f
cc_18 N_VSS_c_15_p N_VDD_c_145_n 3.48826e-19
cc_19 N_VSS_c_7_p N_VDD_c_145_n 0.00955259f
cc_20 N_VSS_c_20_p N_VDD_c_147_n 0.00105775f
cc_21 N_VSS_c_21_p N_VDD_c_148_n 0.00233232f
cc_22 N_VSS_c_4_p N_VDD_c_148_n 9.47758e-19
cc_23 N_VSS_c_13_p N_VDD_c_150_n 3.69367e-19
cc_24 N_VSS_c_21_p N_VDD_c_150_n 0.00161703f
cc_25 N_VSS_c_4_p N_VDD_c_150_n 2.24973e-19
cc_26 N_VSS_c_7_p N_VDD_c_150_n 0.00142089f
cc_27 N_VSS_c_27_p N_VDD_c_150_n 0.00431851f
cc_28 N_VSS_c_28_p N_VDD_c_150_n 7.74609e-19
cc_29 N_VSS_c_3_p N_VDD_c_156_n 0.00179097f
cc_30 N_VSS_c_30_p N_VDD_c_156_n 3.92901e-19
cc_31 N_VSS_c_31_p N_VDD_c_156_n 8.83788e-19
cc_32 N_VSS_c_12_p N_VDD_c_159_n 3.71132e-19
cc_33 N_VSS_c_31_p N_VDD_c_159_n 0.00141228f
cc_34 N_VSS_c_34_p N_VDD_c_159_n 0.00114511f
cc_35 N_VSS_c_35_p N_VDD_c_159_n 0.00431473f
cc_36 N_VSS_c_36_p N_VDD_c_159_n 0.00338293f
cc_37 N_VSS_c_37_p N_VDD_c_159_n 7.74609e-19
cc_38 N_VSS_c_35_p N_VDD_c_165_n 0.00147849f
cc_39 N_VSS_c_21_p N_VDD_c_166_n 9.29349e-19
cc_40 N_VSS_c_4_p N_VDD_c_166_n 3.79458e-19
cc_41 N_VSS_c_41_p N_VDD_c_168_n 2.72411e-19
cc_42 N_VSS_c_42_p N_VDD_c_168_n 3.23198e-19
cc_43 N_VSS_c_27_p N_VDD_c_168_n 0.00448754f
cc_44 N_VSS_c_44_p N_VDD_c_171_n 4.01154e-19
cc_45 N_VSS_c_42_p N_VDD_c_172_n 0.00187494f
cc_46 N_VSS_c_46_p N_VDD_c_172_n 0.00427673f
cc_47 N_VSS_c_47_p N_VDD_c_172_n 0.00924147f
cc_48 N_VSS_c_48_p N_VDD_c_172_n 9.16632e-19
cc_49 N_VSS_c_31_p N_VDD_c_176_n 4.35319e-19
cc_50 N_VSS_c_34_p N_VDD_c_176_n 4.7255e-19
cc_51 N_VSS_c_36_p N_VDD_c_176_n 0.00107125f
cc_52 N_VSS_c_47_p N_VDD_c_176_n 0.00412661f
cc_53 N_VSS_c_3_p N_VDD_c_180_n 6.19689e-19
cc_54 N_VSS_c_54_p N_VDD_c_180_n 3.8721e-19
cc_55 N_VSS_c_15_p N_VDD_c_182_n 0.00178973f
cc_56 N_VSS_c_7_p N_VDD_c_182_n 2.411e-19
cc_57 N_VSS_c_7_p N_VDD_c_184_n 0.00122269f
cc_58 N_VSS_c_27_p N_VDD_c_185_n 0.00106206f
cc_59 N_VSS_c_47_p N_VDD_c_186_n 0.00116512f
cc_60 N_VSS_c_3_p N_VDD_c_187_n 3.86162e-19
cc_61 N_VSS_c_54_p N_VDD_c_187_n 6.0892e-19
cc_62 N_VSS_c_3_p N_VDD_c_189_n 5.2607e-19
cc_63 N_VSS_c_31_p N_VDD_c_189_n 3.48267e-19
cc_64 N_VSS_c_34_p N_VDD_c_189_n 6.489e-19
cc_65 N_VSS_c_21_p N_VDD_c_192_n 3.48267e-19
cc_66 N_VSS_c_4_p N_VDD_c_192_n 6.20986e-19
cc_67 N_VSS_c_14_p N_CKN_c_242_n 3.43419e-19
cc_68 N_VSS_c_15_p N_CKN_c_242_n 3.48267e-19
cc_69 N_VSS_c_15_p N_CKN_c_244_n 0.00109746f
cc_70 N_VSS_c_3_p N_CKN_c_244_n 6.97825e-19
cc_71 N_VSS_c_7_p N_CKN_c_244_n 3.92176e-19
cc_72 N_VSS_c_47_p N_CKN_c_244_n 3.27346e-19
cc_73 N_VSS_c_47_p N_CKN_c_248_n 0.00111539f
cc_74 N_VSS_c_3_p N_CKN_c_249_n 0.00232042f
cc_75 N_VSS_c_30_p N_CKN_c_249_n 5.94801e-19
cc_76 N_VSS_c_31_p N_CKN_c_249_n 3.31491e-19
cc_77 N_VSS_c_7_p N_CKN_c_249_n 0.00107666f
cc_78 N_VSS_c_78_p N_CKN_c_249_n 5.98734e-19
cc_79 N_VSS_c_35_p N_CKN_c_249_n 6.19556e-19
cc_80 N_VSS_c_27_p N_CKN_c_249_n 7.49546e-19
cc_81 N_VSS_c_81_p N_D_c_279_n 5.28294e-19
cc_82 N_VSS_XI13.X0_PGD N_D_c_280_n 3.99797e-19
cc_83 N_VSS_c_3_p N_D_c_281_n 6.13924e-19
cc_84 N_VSS_c_54_p N_D_c_281_n 3.48267e-19
cc_85 N_VSS_c_4_p N_D_c_281_n 2.1322e-19
cc_86 N_VSS_c_3_p N_D_c_284_n 3.48267e-19
cc_87 N_VSS_c_21_p N_D_c_284_n 2.1322e-19
cc_88 N_VSS_c_54_p N_D_c_284_n 6.88619e-19
cc_89 N_VSS_XI5.X0_PGD N_X_c_303_n 4.09718e-19
cc_90 N_VSS_c_41_p N_X_c_304_n 3.43419e-19
cc_91 N_VSS_c_42_p N_X_c_304_n 3.48267e-19
cc_92 N_VSS_c_41_p N_X_c_306_n 3.48267e-19
cc_93 N_VSS_c_3_p N_X_c_306_n 4.71026e-19
cc_94 N_VSS_c_42_p N_X_c_306_n 5.71987e-19
cc_95 N_VSS_c_47_p N_X_c_306_n 3.92273e-19
cc_96 N_VSS_c_3_p N_X_c_310_n 0.00157847f
cc_97 N_VSS_c_47_p N_X_c_310_n 2.88807e-19
cc_98 N_VSS_c_3_p N_X_c_312_n 3.48267e-19
cc_99 N_VSS_c_99_p N_Q_c_349_n 3.43419e-19
cc_100 N_VSS_c_30_p N_Q_c_349_n 3.48267e-19
cc_101 N_VSS_c_30_p Q 5.37696e-19
cc_102 N_CK_c_106_n N_VDD_XI0.X0_PGD 4.20343e-19
cc_103 N_CK_XI13.X0_PGS N_VDD_XI12.X0_PGD 2.44781e-19
cc_104 N_CK_c_107_n N_VDD_c_140_n 2.44781e-19
cc_105 N_CK_c_107_n N_VDD_c_197_n 2.19802e-19
cc_106 CK N_VDD_c_141_n 5.04211e-19
cc_107 N_CK_c_114_p N_VDD_c_141_n 5.29229e-19
cc_108 N_CK_c_106_n N_VDD_c_145_n 0.00150929f
cc_109 CK N_VDD_c_145_n 0.00141439f
cc_110 N_CK_c_114_p N_VDD_c_145_n 0.0012022f
cc_111 N_CK_XI13.X0_PGS N_VDD_c_148_n 2.48209e-19
cc_112 N_CK_c_107_n N_VDD_c_148_n 5.56076e-19
cc_113 CK N_VDD_c_148_n 3.85155e-19
cc_114 N_CK_c_114_p N_VDD_c_148_n 2.72301e-19
cc_115 CK N_VDD_c_180_n 2.86209e-19
cc_116 N_CK_c_114_p N_VDD_c_180_n 2.18105e-19
cc_117 N_CK_c_124_p N_VDD_c_187_n 5.26604e-19
cc_118 CK N_VDD_c_187_n 2.1322e-19
cc_119 N_CK_XI13.X0_PGS N_CKN_XI12.X0_PGS 4.11563e-19
cc_120 N_CK_XI13.X0_PGS N_CKN_c_257_n 2.73384e-19
cc_121 N_CK_c_106_n N_CKN_c_242_n 7.69306e-19
cc_122 N_CK_XI13.X0_PGS N_D_XI13.X0_CG 4.28946e-19
cc_123 N_CK_XI13.X0_PGS N_D_XI12.X0_CG 2.59344e-19
cc_124 N_CK_XI13.X0_PGS N_D_c_284_n 0.00300565f
cc_125 N_CK_XI13.X0_PGS N_X_XI5.X0_CG 2.61247e-19
cc_126 N_CK_XI13.X0_PGS N_X_c_314_n 4.55333e-19
cc_127 N_CK_XI13.X0_PGS N_X_c_312_n 0.00630896f
cc_128 N_VDD_c_172_n N_CKN_XI12.X0_PGS 8.30122e-19
cc_129 N_VDD_c_172_n N_CKN_c_257_n 8.21431e-19
cc_130 N_VDD_c_197_n N_CKN_c_242_n 3.43419e-19
cc_131 N_VDD_c_145_n N_CKN_c_242_n 2.72411e-19
cc_132 N_VDD_c_197_n N_CKN_c_244_n 3.48267e-19
cc_133 N_VDD_c_141_n N_CKN_c_244_n 6.86019e-19
cc_134 N_VDD_c_145_n N_CKN_c_244_n 2.91445e-19
cc_135 N_VDD_c_148_n N_CKN_c_244_n 5.37696e-19
cc_136 N_VDD_c_180_n N_CKN_c_244_n 6.42405e-19
cc_137 N_VDD_c_172_n N_CKN_c_248_n 7.71262e-19
cc_138 N_VDD_c_166_n N_CKN_c_249_n 2.24632e-19
cc_139 N_VDD_XI12.X0_PGD N_D_c_280_n 4.09718e-19
cc_140 N_VDD_XI4.X0_PGD N_X_c_303_n 3.98597e-19
cc_141 N_VDD_c_224_p N_X_c_317_n 4.97416e-19
cc_142 N_VDD_c_197_n N_X_c_304_n 3.43419e-19
cc_143 N_VDD_c_148_n N_X_c_304_n 3.48267e-19
cc_144 N_VDD_c_150_n N_X_c_304_n 2.72411e-19
cc_145 N_VDD_c_197_n N_X_c_306_n 3.48267e-19
cc_146 N_VDD_c_148_n N_X_c_306_n 6.94315e-19
cc_147 N_VDD_c_150_n N_X_c_306_n 3.78778e-19
cc_148 N_VDD_c_172_n N_X_c_306_n 0.00131866f
cc_149 N_VDD_c_156_n N_X_c_310_n 2.90053e-19
cc_150 N_VDD_c_172_n N_X_c_310_n 2.02855e-19
cc_151 N_VDD_c_189_n N_X_c_310_n 2.26379e-19
cc_152 N_VDD_c_156_n N_X_c_312_n 2.28697e-19
cc_153 N_VDD_c_236_p N_Q_c_349_n 3.43419e-19
cc_154 N_VDD_c_159_n N_Q_c_349_n 2.74986e-19
cc_155 N_VDD_c_171_n N_Q_c_349_n 3.72199e-19
cc_156 N_VDD_c_236_p Q 3.48267e-19
cc_157 N_VDD_c_159_n Q 3.66281e-19
cc_158 N_VDD_c_171_n Q 7.06537e-19
cc_159 N_CKN_XI12.X0_PGS N_D_XI12.X0_CG 0.00419505f
cc_160 N_CKN_c_249_n N_D_c_281_n 2.01502e-19
cc_161 N_CKN_XI12.X0_PGS N_X_c_303_n 0.00422719f
cc_162 N_CKN_c_257_n N_X_c_330_n 5.71169e-19
cc_163 N_CKN_c_249_n N_X_c_330_n 0.00194262f
cc_164 N_CKN_c_244_n N_X_c_306_n 7.35688e-19
cc_165 N_CKN_c_248_n N_X_c_306_n 8.08281e-19
cc_166 N_CKN_c_249_n N_X_c_306_n 7.34542e-19
cc_167 N_CKN_c_249_n N_X_c_310_n 8.56658e-19
cc_168 N_D_c_280_n N_X_c_303_n 0.00477695f
cc_169 N_D_c_280_n N_X_c_304_n 6.90199e-19
cc_170 N_D_c_280_n N_X_c_330_n 4.21501e-19
cc_171 N_D_c_280_n N_X_c_306_n 3.40033e-19
cc_172 N_D_c_281_n N_X_c_306_n 0.00151909f
cc_173 N_D_c_284_n N_X_c_306_n 0.00104518f
cc_174 N_D_c_281_n N_X_c_310_n 0.00146206f
cc_175 N_D_c_284_n N_X_c_310_n 0.00103457f
cc_176 N_D_c_281_n N_X_c_312_n 4.56568e-19
cc_177 N_D_c_284_n N_X_c_312_n 0.00383269f
cc_178 N_X_c_303_n N_Q_c_349_n 6.90199e-19
cc_179 N_X_c_330_n N_Q_c_349_n 3.5757e-19
cc_180 N_X_c_330_n Q 5.52904e-19
*
.ends
*
*
.subckt DFFQ1_HPNW12 CK D Q VDD VSS
xgate (VSS CK VDD D Q) G3_DFFQ1_N3
.ends
*
* File: G1_INV1_N3.pex.netlist
* Created: Fri Feb 25 16:26:51 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G1_INV1_N3_VDD 2 5 15 23 28 30 34 37 43 Vss
c22 43 Vss 0.00440656f
c23 34 Vss 7.98732e-19
c24 30 Vss 0.00491201f
c25 28 Vss 0.0026398f
c26 26 Vss 0.00168274f
c27 23 Vss 0.00814922f
c28 15 Vss 0.0356247f
c29 14 Vss 0.102427f
c30 5 Vss 0.382574f
r31 34 43 1.16709
r32 32 34 2.41736
r33 31 37 0.326018
r34 30 32 0.652036
r35 30 31 7.46046
r36 26 37 0.326018
r37 26 28 6.4185
r38 23 28 1.16709
r39 17 43 0.0476429
r40 15 17 1.45875
r41 14 18 0.652036
r42 14 17 1.45875
r43 11 15 0.652036
r44 5 18 5.1348
r45 5 11 5.1348
r46 2 23 0.123773
.ends

.subckt PM_G1_INV1_N3_A 2 4 12 24 27 Vss
c6 27 Vss 0.00733896f
c7 24 Vss 1.81646e-19
c8 12 Vss 0.229828f
c9 9 Vss 0.180667f
c10 7 Vss 0.0247918f
c11 4 Vss 0.193588f
r12 24 27 1.16709
r13 15 27 0.0476429
r14 13 15 0.326018
r15 13 15 0.1167
r16 12 16 0.652036
r17 12 15 6.7686
r18 9 27 0.357321
r19 7 15 0.326018
r20 7 9 0.40845
r21 4 16 5.1348
r22 2 9 4.72635
.ends

.subckt PM_G1_INV1_N3_VSS 3 6 14 24 27 32 37 49 50 56 Vss
c23 51 Vss 0.0012698f
c24 50 Vss 6.56512e-19
c25 49 Vss 0.00353949f
c26 37 Vss 0.00390919f
c27 32 Vss 0.00198602f
c28 27 Vss 8.43451e-19
c29 24 Vss 0.0100686f
c30 15 Vss 0.0359156f
c31 14 Vss 0.0994171f
c32 3 Vss 0.381612f
r33 51 56 0.326018
r34 49 56 0.326018
r35 49 50 7.46046
r36 45 50 0.652036
r37 32 51 6.4185
r38 27 37 1.16709
r39 27 45 2.41736
r40 24 32 1.16709
r41 17 37 0.0476429
r42 15 17 1.45875
r43 14 18 0.652036
r44 14 17 1.45875
r45 11 15 0.652036
r46 6 24 0.123773
r47 3 18 5.1348
r48 3 11 5.1348
.ends

.subckt PM_G1_INV1_N3_Z 2 4 13 19 Vss
c11 13 Vss 0.00499164f
c12 4 Vss 0.00143493f
r13 16 19 0.0364688
r14 13 16 1.16709
r15 4 13 0.123773
r16 2 13 0.123773
.ends

.subckt G1_INV1_N3  VDD A VSS Z
*
* Z	Z
* VSS	VSS
* A	A
* VDD	VDD
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_A_XI6.X0_CG N_VSS_XI6.X0_PGD
+ N_VDD_XI6.X0_S TIGFET_HPNW12
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_A_XI5.X0_CG N_VDD_XI5.X0_PGD
+ N_VSS_XI5.X0_S TIGFET_HPNW12
*
x_PM_G1_INV1_N3_VDD N_VDD_XI6.X0_S N_VDD_XI5.X0_PGD N_VDD_c_4_p N_VDD_c_17_p
+ N_VDD_c_3_p N_VDD_c_5_p N_VDD_c_8_p VDD N_VDD_c_9_p Vss PM_G1_INV1_N3_VDD
x_PM_G1_INV1_N3_A N_A_XI6.X0_CG N_A_XI5.X0_CG N_A_c_23_n A N_A_c_26_p Vss
+ PM_G1_INV1_N3_A
x_PM_G1_INV1_N3_VSS N_VSS_XI6.X0_PGD N_VSS_XI5.X0_S N_VSS_c_31_n N_VSS_c_48_p
+ N_VSS_c_33_n N_VSS_c_37_n N_VSS_c_39_n N_VSS_c_42_n N_VSS_c_43_n VSS Vss
+ PM_G1_INV1_N3_VSS
x_PM_G1_INV1_N3_Z N_Z_XI6.X0_D N_Z_XI5.X0_D N_Z_c_52_n Z Vss PM_G1_INV1_N3_Z
cc_1 N_VDD_XI5.X0_PGD N_A_c_23_n 4.31283e-19
cc_2 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.00199939f
cc_3 N_VDD_c_3_p N_VSS_XI6.X0_PGD 4.23795e-19
cc_4 N_VDD_c_4_p N_VSS_c_31_n 0.00199939f
cc_5 N_VDD_c_5_p N_VSS_c_31_n 5.08727e-19
cc_6 N_VDD_c_3_p N_VSS_c_33_n 0.00302944f
cc_7 N_VDD_c_5_p N_VSS_c_33_n 0.00141897f
cc_8 N_VDD_c_8_p N_VSS_c_33_n 9.31072e-19
cc_9 N_VDD_c_9_p N_VSS_c_33_n 3.48267e-19
cc_10 N_VDD_c_3_p N_VSS_c_37_n 7.58061e-19
cc_11 N_VDD_c_8_p N_VSS_c_37_n 0.00105766f
cc_12 N_VDD_c_3_p N_VSS_c_39_n 9.55109e-19
cc_13 N_VDD_c_5_p N_VSS_c_39_n 0.00103739f
cc_14 N_VDD_c_9_p N_VSS_c_39_n 6.46219e-19
cc_15 N_VDD_c_5_p N_VSS_c_42_n 0.0059288f
cc_16 N_VDD_c_5_p N_VSS_c_43_n 0.00172731f
cc_17 N_VDD_c_17_p N_Z_c_52_n 3.43419e-19
cc_18 N_VDD_c_3_p N_Z_c_52_n 3.48267e-19
cc_19 N_VDD_c_5_p N_Z_c_52_n 2.60012e-19
cc_20 N_VDD_c_17_p Z 3.48267e-19
cc_21 N_VDD_c_3_p Z 7.09569e-19
cc_22 N_VDD_c_5_p Z 3.45966e-19
cc_23 N_A_c_23_n N_VSS_XI6.X0_PGD 4.31283e-19
cc_24 A N_VSS_c_33_n 3.42414e-19
cc_25 N_A_c_26_p N_VSS_c_33_n 2.30774e-19
cc_26 A N_VSS_c_39_n 2.30774e-19
cc_27 N_A_c_23_n N_Z_c_52_n 7.69306e-19
cc_28 N_VSS_c_48_p N_Z_c_52_n 3.43419e-19
cc_29 N_VSS_c_37_n N_Z_c_52_n 3.48267e-19
cc_30 N_VSS_c_37_n Z 8.23589e-19
cc_31 N_VSS_c_42_n Z 2.18525e-19
*
.ends
*
*
.subckt INV1_HPNW12 A Y VDD VSS
xgate (VDD A VSS Y) G1_INV1_N3
.ends
*
* File: G3_LATQ1_N3.pex.netlist
* Created: Tue Apr  5 12:00:00 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_LATQ1_N3_VDD 2 4 6 8 10 12 14 16 31 42 48 58 63 66 68 69 70 71 72
+ 75 77 81 85 90 92 98 103 Vss
c82 103 Vss 0.00476181f
c83 98 Vss 0.00486653f
c84 90 Vss 2.39889e-19
c85 85 Vss 0.00253232f
c86 83 Vss 0.0017055f
c87 81 Vss 0.00108379f
c88 77 Vss 0.0043713f
c89 75 Vss 8.9379e-19
c90 72 Vss 8.65746e-19
c91 71 Vss 0.00223415f
c92 70 Vss 8.64769e-19
c93 69 Vss 0.00576876f
c94 68 Vss 0.0113641f
c95 66 Vss 0.00582672f
c96 63 Vss 0.00607435f
c97 58 Vss 0.00819566f
c98 53 Vss 0.0307825f
c99 48 Vss 0.230506f
c100 44 Vss 1.68267e-19
c101 42 Vss 0.0357228f
c102 41 Vss 0.0656875f
c103 32 Vss 0.0359366f
c104 31 Vss 0.101312f
c105 16 Vss 0.00143493f
c106 14 Vss 0.191707f
c107 10 Vss 0.191287f
c108 8 Vss 0.189707f
c109 6 Vss 0.190072f
c110 4 Vss 0.189718f
r111 83 92 0.326018
r112 83 85 6.16843
r113 81 103 1.16709
r114 79 81 2.16729
r115 78 90 0.494161
r116 77 92 0.326018
r117 77 78 7.46046
r118 75 98 1.16709
r119 73 90 0.128424
r120 73 75 2.16729
r121 71 90 0.494161
r122 71 72 4.37625
r123 69 79 0.652036
r124 69 70 10.1279
r125 68 72 0.652036
r126 67 68 18.2969
r127 66 89 2.334
r128 66 67 0.14525
r129 65 70 0.652036
r130 65 66 5.54325
r131 63 85 1.16709
r132 58 89 1.16709
r133 49 53 0.494161
r134 48 50 0.652036
r135 48 49 6.8853
r136 45 53 0.128424
r137 44 103 0.0476429
r138 42 44 1.45875
r139 41 53 0.494161
r140 41 44 1.45875
r141 38 42 0.652036
r142 34 98 0.0476429
r143 32 34 1.45875
r144 31 35 0.652036
r145 31 34 1.45875
r146 28 32 0.652036
r147 16 63 0.123773
r148 14 50 5.1348
r149 12 63 0.123773
r150 10 45 5.1348
r151 8 38 5.1348
r152 6 28 5.1348
r153 4 35 5.1348
r154 2 58 0.123773
.ends

.subckt PM_G3_LATQ1_N3_VSS 2 4 6 8 10 12 14 16 31 32 34 42 48 58 63 66 71 76 81
+ 90 95 104 106 107 108 113 114 119 129 130 132 Vss
c74 130 Vss 3.75522e-19
c75 129 Vss 4.28045e-19
c76 125 Vss 0.00128551f
c77 119 Vss 0.00327372f
c78 114 Vss 8.25631e-19
c79 113 Vss 0.00434469f
c80 108 Vss 8.30816e-19
c81 107 Vss 0.00172205f
c82 106 Vss 0.00206535f
c83 104 Vss 0.00621153f
c84 95 Vss 0.00443295f
c85 90 Vss 0.0041985f
c86 81 Vss 0.00249073f
c87 76 Vss 9.5519e-19
c88 71 Vss 6.07136e-19
c89 66 Vss 0.0013933f
c90 63 Vss 0.0060193f
c91 58 Vss 0.00814768f
c92 53 Vss 0.0307825f
c93 48 Vss 0.231473f
c94 42 Vss 0.0348714f
c95 41 Vss 0.0647879f
c96 34 Vss 8.95828e-20
c97 32 Vss 0.0350852f
c98 31 Vss 0.0994129f
c99 16 Vss 0.191895f
c100 14 Vss 0.00143493f
c101 12 Vss 0.19162f
c102 10 Vss 0.189706f
c103 4 Vss 0.190073f
c104 2 Vss 0.18972f
r105 125 132 0.326018
r106 120 130 0.494161
r107 119 132 0.326018
r108 119 120 7.46046
r109 115 130 0.128424
r110 113 121 0.652036
r111 113 114 10.1279
r112 109 129 0.0828784
r113 107 130 0.494161
r114 107 108 4.37625
r115 106 114 0.652036
r116 105 129 0.551426
r117 105 106 5.50157
r118 104 129 0.551426
r119 103 108 0.652036
r120 103 104 18.3386
r121 81 125 6.16843
r122 76 95 1.16709
r123 76 121 2.16729
r124 71 90 1.16709
r125 71 115 2.16729
r126 66 109 1.82344
r127 63 81 1.16709
r128 58 66 1.16709
r129 49 53 0.494161
r130 48 50 0.652036
r131 48 49 6.8853
r132 45 53 0.128424
r133 44 95 0.0476429
r134 42 44 1.45875
r135 41 53 0.494161
r136 41 44 1.45875
r137 38 42 0.652036
r138 34 90 0.0476429
r139 32 34 1.45875
r140 31 35 0.652036
r141 31 34 1.45875
r142 28 32 0.652036
r143 16 50 5.1348
r144 14 63 0.123773
r145 12 45 5.1348
r146 10 38 5.1348
r147 8 63 0.123773
r148 6 58 0.123773
r149 4 28 5.1348
r150 2 35 5.1348
.ends

.subckt PM_G3_LATQ1_N3_G 2 4 6 14 15 22 31 37 Vss
c24 37 Vss 0.00266632f
c25 31 Vss 6.62558e-19
c26 29 Vss 0.0295325f
c27 22 Vss 0.152777f
c28 15 Vss 0.179526f
c29 14 Vss 2.0264e-19
c30 10 Vss 0.0247918f
c31 6 Vss 0.192371f
c32 4 Vss 0.193138f
c33 2 Vss 0.180487f
r34 34 37 1.16709
r35 31 34 0.0833571
r36 23 29 0.494161
r37 22 24 0.652036
r38 22 23 4.84305
r39 19 29 0.128424
r40 18 37 0.0476429
r41 16 18 0.326018
r42 16 18 0.1167
r43 15 29 0.494161
r44 15 18 6.7686
r45 14 37 0.357321
r46 10 18 0.326018
r47 10 14 0.40845
r48 6 24 5.1348
r49 4 19 5.1348
r50 2 14 4.72635
.ends

.subckt PM_G3_LATQ1_N3_QN 2 4 6 8 20 23 33 37 40 45 48 53 69 Vss
c43 69 Vss 4.86032e-19
c44 53 Vss 0.00238508f
c45 48 Vss 0.00856405f
c46 45 Vss 0.00518251f
c47 40 Vss 0.00103774f
c48 37 Vss 0.0113402f
c49 33 Vss 0.0113402f
c50 23 Vss 2.25442e-19
c51 20 Vss 0.214677f
c52 17 Vss 0.180502f
c53 15 Vss 0.0247918f
c54 4 Vss 0.191818f
r55 65 69 0.652036
r56 48 69 13.7956
r57 48 50 6.4185
r58 45 48 6.4185
r59 40 53 1.16709
r60 40 65 1.83386
r61 37 50 1.16709
r62 33 45 1.16709
r63 23 53 0.0476429
r64 21 23 0.326018
r65 21 23 0.1167
r66 20 24 0.652036
r67 20 23 6.7686
r68 17 53 0.357321
r69 15 23 0.326018
r70 15 17 0.40845
r71 8 37 0.123773
r72 6 33 0.123773
r73 4 24 5.1348
r74 2 17 4.72635
.ends

.subckt PM_G3_LATQ1_N3_GN 2 4 6 12 23 27 29 30 32 39 Vss
c39 39 Vss 0.00500045f
c40 32 Vss 6.08951e-19
c41 30 Vss 6.08791e-19
c42 29 Vss 0.00111596f
c43 27 Vss 0.00109183f
c44 23 Vss 0.00525048f
c45 14 Vss 1.82689e-19
c46 12 Vss 0.163012f
c47 6 Vss 0.285833f
c48 4 Vss 0.00143493f
r49 32 39 1.16709
r50 29 32 0.531835
r51 29 30 1.70882
r52 25 30 0.652036
r53 25 27 5.835
r54 23 27 1.16709
r55 14 39 0.197068
r56 12 16 0.652036
r57 12 14 4.668
r58 6 16 8.4024
r59 4 23 0.123773
r60 2 23 0.123773
.ends

.subckt PM_G3_LATQ1_N3_Q 2 4 13 18 Vss
c12 18 Vss 3.21524e-19
c13 13 Vss 0.00454527f
c14 4 Vss 0.00143493f
r15 13 18 1.16709
r16 4 13 0.123773
r17 2 13 0.123773
.ends

.subckt PM_G3_LATQ1_N3_D 2 4 10 14 Vss
c14 14 Vss 4.85129e-19
c15 10 Vss 1.35847e-19
c16 2 Vss 0.58413f
r17 14 17 0.0416786
r18 10 17 1.16709
r19 4 10 8.9859
r20 2 10 8.9859
.ends

.subckt G3_LATQ1_N3  VDD VSS G Q D
*
* D	D
* Q	Q
* G	G
* VSS	VSS
* VDD	VDD
XI3.X0 N_GN_XI3.X0_D N_VSS_XI3.X0_PGD N_G_XI3.X0_CG N_VSS_XI3.X0_PGS
+ N_VDD_XI3.X0_S TIGFET_HPNW12
XI0.X0 N_Q_XI0.X0_D N_VDD_XI0.X0_PGD N_QN_XI0.X0_CG N_VDD_XI0.X0_PGS
+ N_VSS_XI0.X0_S TIGFET_HPNW12
XI1.X0 N_GN_XI1.X0_D N_VDD_XI1.X0_PGD N_G_XI1.X0_CG N_VDD_XI1.X0_PGS
+ N_VSS_XI1.X0_S TIGFET_HPNW12
XI4.X0 N_Q_XI4.X0_D N_VSS_XI4.X0_PGD N_QN_XI4.X0_CG N_VSS_XI4.X0_PGS
+ N_VDD_XI4.X0_S TIGFET_HPNW12
XI2.X0 N_QN_XI2.X0_D N_VDD_XI2.X0_PGD N_D_XI2.X0_CG N_G_XI2.X0_PGS
+ N_VSS_XI2.X0_S TIGFET_HPNW12
XI5.X0 N_QN_XI5.X0_D N_VSS_XI5.X0_PGD N_D_XI5.X0_CG N_GN_XI5.X0_PGS
+ N_VDD_XI5.X0_S TIGFET_HPNW12
*
x_PM_G3_LATQ1_N3_VDD N_VDD_XI3.X0_S N_VDD_XI0.X0_PGD N_VDD_XI0.X0_PGS
+ N_VDD_XI1.X0_PGD N_VDD_XI1.X0_PGS N_VDD_XI4.X0_S N_VDD_XI2.X0_PGD
+ N_VDD_XI5.X0_S N_VDD_c_9_p N_VDD_c_5_p N_VDD_c_14_p N_VDD_c_69_p N_VDD_c_11_p
+ N_VDD_c_7_p N_VDD_c_13_p N_VDD_c_6_p N_VDD_c_41_p N_VDD_c_18_p N_VDD_c_45_p
+ N_VDD_c_23_p N_VDD_c_10_p N_VDD_c_21_p N_VDD_c_12_p N_VDD_c_44_p VDD
+ N_VDD_c_26_p N_VDD_c_22_p Vss PM_G3_LATQ1_N3_VDD
x_PM_G3_LATQ1_N3_VSS N_VSS_XI3.X0_PGD N_VSS_XI3.X0_PGS N_VSS_XI0.X0_S
+ N_VSS_XI1.X0_S N_VSS_XI4.X0_PGD N_VSS_XI4.X0_PGS N_VSS_XI2.X0_S
+ N_VSS_XI5.X0_PGD N_VSS_c_87_n N_VSS_c_89_n N_VSS_c_131_p N_VSS_c_91_n
+ N_VSS_c_93_n N_VSS_c_95_n N_VSS_c_96_n N_VSS_c_98_n N_VSS_c_101_n
+ N_VSS_c_105_n N_VSS_c_109_n N_VSS_c_111_n N_VSS_c_115_n N_VSS_c_119_n
+ N_VSS_c_121_n N_VSS_c_122_n N_VSS_c_123_n N_VSS_c_124_n N_VSS_c_127_n
+ N_VSS_c_128_n N_VSS_c_129_n N_VSS_c_130_n VSS Vss PM_G3_LATQ1_N3_VSS
x_PM_G3_LATQ1_N3_G N_G_XI3.X0_CG N_G_XI1.X0_CG N_G_XI2.X0_PGS N_G_c_162_n
+ N_G_c_158_n N_G_c_159_n G N_G_c_161_n Vss PM_G3_LATQ1_N3_G
x_PM_G3_LATQ1_N3_QN N_QN_XI0.X0_CG N_QN_XI4.X0_CG N_QN_XI2.X0_D N_QN_XI5.X0_D
+ N_QN_c_181_n N_QN_c_182_n N_QN_c_196_n N_QN_c_183_n N_QN_c_185_n N_QN_c_187_n
+ N_QN_c_189_n N_QN_c_192_n N_QN_c_194_n Vss PM_G3_LATQ1_N3_QN
x_PM_G3_LATQ1_N3_GN N_GN_XI3.X0_D N_GN_XI1.X0_D N_GN_XI5.X0_PGS N_GN_c_224_n
+ N_GN_c_225_n N_GN_c_228_n N_GN_c_244_n N_GN_c_250_n N_GN_c_252_n N_GN_c_245_n
+ Vss PM_G3_LATQ1_N3_GN
x_PM_G3_LATQ1_N3_Q N_Q_XI0.X0_D N_Q_XI4.X0_D N_Q_c_263_n Q Vss PM_G3_LATQ1_N3_Q
x_PM_G3_LATQ1_N3_D N_D_XI2.X0_CG N_D_XI5.X0_CG N_D_c_280_n D Vss
+ PM_G3_LATQ1_N3_D
cc_1 N_VDD_XI1.X0_PGD N_VSS_XI3.X0_PGD 0.00203852f
cc_2 N_VDD_XI0.X0_PGS N_VSS_XI3.X0_PGS 2.44446e-19
cc_3 N_VDD_XI0.X0_PGD N_VSS_XI4.X0_PGD 0.00203076f
cc_4 N_VDD_XI2.X0_PGD N_VSS_XI5.X0_PGD 2.44446e-19
cc_5 N_VDD_c_5_p N_VSS_c_87_n 0.00203852f
cc_6 N_VDD_c_6_p N_VSS_c_87_n 3.89167e-19
cc_7 N_VDD_c_7_p N_VSS_c_89_n 3.80615e-19
cc_8 N_VDD_c_6_p N_VSS_c_89_n 3.89167e-19
cc_9 N_VDD_c_9_p N_VSS_c_91_n 0.00203076f
cc_10 N_VDD_c_10_p N_VSS_c_91_n 3.00073e-19
cc_11 N_VDD_c_11_p N_VSS_c_93_n 2.19802e-19
cc_12 N_VDD_c_12_p N_VSS_c_93_n 8.58125e-19
cc_13 N_VDD_c_13_p N_VSS_c_95_n 9.5668e-19
cc_14 N_VDD_c_14_p N_VSS_c_96_n 2.19802e-19
cc_15 N_VDD_c_11_p N_VSS_c_96_n 2.80254e-19
cc_16 N_VDD_c_7_p N_VSS_c_98_n 4.06916e-19
cc_17 N_VDD_c_13_p N_VSS_c_98_n 0.00165395f
cc_18 N_VDD_c_18_p N_VSS_c_98_n 3.5277e-19
cc_19 N_VDD_c_7_p N_VSS_c_101_n 9.31121e-19
cc_20 N_VDD_c_6_p N_VSS_c_101_n 0.00161703f
cc_21 N_VDD_c_21_p N_VSS_c_101_n 7.09654e-19
cc_22 N_VDD_c_22_p N_VSS_c_101_n 3.48267e-19
cc_23 N_VDD_c_23_p N_VSS_c_105_n 9.52068e-19
cc_24 N_VDD_c_10_p N_VSS_c_105_n 0.00141228f
cc_25 N_VDD_c_12_p N_VSS_c_105_n 0.00257912f
cc_26 N_VDD_c_26_p N_VSS_c_105_n 3.48267e-19
cc_27 N_VDD_c_7_p N_VSS_c_109_n 3.32876e-19
cc_28 N_VDD_c_21_p N_VSS_c_109_n 8.43845e-19
cc_29 N_VDD_c_7_p N_VSS_c_111_n 4.24454e-19
cc_30 N_VDD_c_6_p N_VSS_c_111_n 2.26455e-19
cc_31 N_VDD_c_21_p N_VSS_c_111_n 3.84769e-19
cc_32 N_VDD_c_22_p N_VSS_c_111_n 6.489e-19
cc_33 N_VDD_c_23_p N_VSS_c_115_n 3.82294e-19
cc_34 N_VDD_c_10_p N_VSS_c_115_n 0.00114511f
cc_35 N_VDD_c_12_p N_VSS_c_115_n 9.55109e-19
cc_36 N_VDD_c_26_p N_VSS_c_115_n 6.46219e-19
cc_37 N_VDD_c_7_p N_VSS_c_119_n 0.00540208f
cc_38 N_VDD_c_13_p N_VSS_c_119_n 0.00786235f
cc_39 N_VDD_c_13_p N_VSS_c_121_n 0.00445899f
cc_40 N_VDD_c_6_p N_VSS_c_122_n 0.00348718f
cc_41 N_VDD_c_41_p N_VSS_c_123_n 0.00106807f
cc_42 N_VDD_c_18_p N_VSS_c_124_n 0.00356332f
cc_43 N_VDD_c_10_p N_VSS_c_124_n 0.00600653f
cc_44 N_VDD_c_44_p N_VSS_c_124_n 0.00103147f
cc_45 N_VDD_c_45_p N_VSS_c_127_n 0.00106428f
cc_46 N_VDD_c_6_p N_VSS_c_128_n 0.00586992f
cc_47 N_VDD_c_13_p N_VSS_c_129_n 9.16632e-19
cc_48 N_VDD_c_6_p N_VSS_c_130_n 7.74609e-19
cc_49 N_VDD_c_14_p N_G_XI2.X0_PGS 0.00172513f
cc_50 N_VDD_XI1.X0_PGD N_G_c_158_n 3.99191e-19
cc_51 N_VDD_XI1.X0_PGS N_G_c_159_n 4.09718e-19
cc_52 N_VDD_c_13_p G 5.04211e-19
cc_53 N_VDD_c_13_p N_G_c_161_n 5.56409e-19
cc_54 N_VDD_XI0.X0_PGD N_QN_c_181_n 4.09718e-19
cc_55 N_VDD_c_26_p N_QN_c_182_n 6.34963e-19
cc_56 N_VDD_c_11_p N_QN_c_183_n 3.43419e-19
cc_57 N_VDD_c_12_p N_QN_c_183_n 3.48267e-19
cc_58 N_VDD_c_13_p N_QN_c_185_n 4.49462e-19
cc_59 N_VDD_c_26_p N_QN_c_185_n 2.10618e-19
cc_60 N_VDD_c_11_p N_QN_c_187_n 3.48267e-19
cc_61 N_VDD_c_12_p N_QN_c_187_n 9.04108e-19
cc_62 N_VDD_c_6_p N_QN_c_189_n 3.28643e-19
cc_63 N_VDD_c_10_p N_QN_c_189_n 2.94643e-19
cc_64 N_VDD_c_12_p N_QN_c_189_n 3.47038e-19
cc_65 N_VDD_c_13_p N_QN_c_192_n 2.92308e-19
cc_66 N_VDD_c_23_p N_QN_c_192_n 2.28697e-19
cc_67 N_VDD_c_13_p N_QN_c_194_n 3.90734e-19
cc_68 N_VDD_c_11_p N_GN_c_224_n 3.11705e-19
cc_69 N_VDD_c_69_p N_GN_c_225_n 3.43419e-19
cc_70 N_VDD_c_7_p N_GN_c_225_n 3.72199e-19
cc_71 N_VDD_c_6_p N_GN_c_225_n 2.74986e-19
cc_72 N_VDD_c_69_p N_GN_c_228_n 3.48267e-19
cc_73 N_VDD_c_7_p N_GN_c_228_n 7.94301e-19
cc_74 N_VDD_c_13_p N_GN_c_228_n 0.00122181f
cc_75 N_VDD_c_6_p N_GN_c_228_n 3.82604e-19
cc_76 N_VDD_c_11_p N_Q_c_263_n 3.43419e-19
cc_77 N_VDD_c_10_p N_Q_c_263_n 2.74986e-19
cc_78 N_VDD_c_12_p N_Q_c_263_n 3.48267e-19
cc_79 N_VDD_c_11_p Q 3.48267e-19
cc_80 N_VDD_c_10_p Q 3.66281e-19
cc_81 N_VDD_c_12_p Q 7.09569e-19
cc_82 N_VDD_c_14_p N_D_XI2.X0_CG 4.32953e-19
cc_83 N_VSS_c_131_p N_G_c_162_n 5.35095e-19
cc_84 N_VSS_XI3.X0_PGD N_G_c_158_n 4.09718e-19
cc_85 N_VSS_c_111_n G 2.15082e-19
cc_86 N_VSS_c_119_n G 2.86445e-19
cc_87 N_VSS_c_101_n N_G_c_161_n 2.15082e-19
cc_88 N_VSS_XI4.X0_PGD N_QN_c_181_n 3.99191e-19
cc_89 N_VSS_c_96_n N_QN_c_196_n 3.43419e-19
cc_90 N_VSS_c_109_n N_QN_c_196_n 3.48267e-19
cc_91 N_VSS_c_96_n N_QN_c_187_n 3.48267e-19
cc_92 N_VSS_c_109_n N_QN_c_187_n 8.62542e-19
cc_93 N_VSS_c_109_n N_QN_c_189_n 5.58212e-19
cc_94 N_VSS_c_124_n N_QN_c_189_n 4.58442e-19
cc_95 N_VSS_c_128_n N_QN_c_189_n 6.13056e-19
cc_96 N_VSS_c_101_n N_QN_c_194_n 3.59967e-19
cc_97 N_VSS_c_119_n N_QN_c_194_n 0.00182171f
cc_98 N_VSS_c_93_n N_GN_XI5.X0_PGS 0.00172853f
cc_99 N_VSS_XI4.X0_PGS N_GN_c_224_n 6.66551e-19
cc_100 N_VSS_c_96_n N_GN_c_225_n 3.43419e-19
cc_101 N_VSS_c_109_n N_GN_c_225_n 3.48267e-19
cc_102 N_VSS_c_96_n N_GN_c_228_n 3.48267e-19
cc_103 N_VSS_c_109_n N_GN_c_228_n 4.99861e-19
cc_104 N_VSS_c_119_n N_GN_c_228_n 7.12611e-19
cc_105 N_VSS_c_95_n N_Q_c_263_n 3.43419e-19
cc_106 N_VSS_c_98_n N_Q_c_263_n 3.48267e-19
cc_107 N_VSS_c_98_n Q 8.15956e-19
cc_108 N_VSS_c_93_n N_D_XI2.X0_CG 4.32953e-19
cc_109 N_G_c_158_n N_QN_c_181_n 0.00400131f
cc_110 G N_QN_c_185_n 4.48861e-19
cc_111 N_G_c_161_n N_QN_c_185_n 4.54925e-19
cc_112 G N_QN_c_192_n 4.56568e-19
cc_113 N_G_c_161_n N_QN_c_192_n 0.00268575f
cc_114 N_G_c_159_n N_GN_c_224_n 0.00878732f
cc_115 N_G_c_158_n N_GN_c_225_n 6.90199e-19
cc_116 N_G_c_158_n N_GN_c_228_n 3.82175e-19
cc_117 G N_GN_c_228_n 0.00151253f
cc_118 N_G_c_161_n N_GN_c_228_n 9.72448e-19
cc_119 N_G_c_158_n N_GN_c_244_n 4.1347e-19
cc_120 N_G_c_158_n N_GN_c_245_n 0.00397074f
cc_121 N_G_c_161_n N_GN_c_245_n 2.41671e-19
cc_122 N_G_XI2.X0_PGS N_D_XI2.X0_CG 0.00435077f
cc_123 N_QN_c_181_n N_GN_XI5.X0_PGS 0.00196434f
cc_124 N_QN_c_187_n N_GN_c_228_n 0.00124016f
cc_125 N_QN_c_189_n N_GN_c_244_n 0.00100851f
cc_126 N_QN_c_181_n N_GN_c_250_n 4.04137e-19
cc_127 N_QN_c_189_n N_GN_c_250_n 0.00133182f
cc_128 N_QN_c_189_n N_GN_c_252_n 0.00102929f
cc_129 N_QN_c_181_n N_GN_c_245_n 0.00341994f
cc_130 N_QN_c_192_n N_GN_c_245_n 2.75519e-19
cc_131 N_QN_c_181_n N_Q_c_263_n 6.90199e-19
cc_132 N_QN_c_181_n N_D_XI2.X0_CG 3.26559e-19
cc_133 N_QN_c_187_n N_D_XI2.X0_CG 0.0010503f
cc_134 N_QN_c_187_n N_D_c_280_n 0.00130556f
cc_135 N_QN_c_187_n D 0.00141415f
cc_136 N_QN_c_189_n D 0.00146947f
cc_137 N_GN_c_250_n N_Q_c_263_n 3.29741e-19
cc_138 N_GN_c_250_n Q 3.9897e-19
cc_139 N_GN_XI5.X0_PGS N_D_XI2.X0_CG 0.0048787f
cc_140 N_GN_c_224_n N_D_c_280_n 0.00333193f
cc_141 N_GN_c_252_n N_D_c_280_n 3.73302e-19
cc_142 N_GN_c_245_n N_D_c_280_n 8.5422e-19
cc_143 N_GN_c_252_n D 2.85187e-19
cc_144 N_GN_c_245_n D 3.48267e-19
*
.ends
*
*
.subckt LATQ1_HPNW12 D G Q VDD VSS
xgate (VDD VSS G Q D) G3_LATQ1_N3
.ends
*
* File: G4_MAJ3_N3.pex.netlist
* Created: Fri Mar  4 11:51:04 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MAJ3_N3_VDD 2 4 7 11 27 28 30 31 32 44 48 52 54 56 57 58 61 65 67
+ 69 70 73 77 79 80 90 95 Vss
c76 95 Vss 0.00472824f
c77 90 Vss 0.00466016f
c78 80 Vss 4.52364e-19
c79 79 Vss 4.28405e-19
c80 77 Vss 4.68316e-19
c81 73 Vss 0.00105057f
c82 70 Vss 8.64769e-19
c83 69 Vss 0.00576436f
c84 67 Vss 0.00145931f
c85 61 Vss 0.00146297f
c86 58 Vss 8.64769e-19
c87 57 Vss 0.00590519f
c88 56 Vss 0.0027558f
c89 54 Vss 0.0069447f
c90 52 Vss 0.00282697f
c91 48 Vss 0.00810125f
c92 44 Vss 0.0099068f
c93 32 Vss 0.0356247f
c94 31 Vss 0.10084f
c95 28 Vss 0.0356247f
c96 27 Vss 0.100978f
c97 11 Vss 0.376343f
c98 7 Vss 0.374237f
r99 77 95 1.16709
r100 75 77 2.16729
r101 73 90 1.16709
r102 71 73 2.16729
r103 69 75 0.652036
r104 69 70 10.1279
r105 65 67 1.167
r106 63 80 0.0828784
r107 63 65 0.656438
r108 59 79 0.0828784
r109 59 61 1.82344
r110 57 71 0.652036
r111 57 58 10.1279
r112 56 70 0.652036
r113 55 80 0.551426
r114 55 56 5.50157
r115 54 80 0.551426
r116 53 79 0.551426
r117 53 54 11.5033
r118 52 79 0.551426
r119 51 58 0.652036
r120 51 52 5.50157
r121 48 67 1.16709
r122 44 61 1.16709
r123 34 95 0.0476429
r124 32 34 1.45875
r125 31 38 0.652036
r126 31 34 1.45875
r127 30 90 0.0476429
r128 28 30 1.45875
r129 27 35 0.652036
r130 27 30 1.45875
r131 24 32 0.652036
r132 21 28 0.652036
r133 11 38 5.1348
r134 11 24 5.1348
r135 7 35 5.1348
r136 7 21 5.1348
r137 4 48 0.123773
r138 2 44 0.123773
.ends

.subckt PM_G4_MAJ3_N3_VSS 3 7 10 12 27 28 31 32 45 49 52 57 62 67 70 73 78 91 92
+ 93 94 95 104 114 115 117 Vss
c81 115 Vss 3.75522e-19
c82 114 Vss 3.75522e-19
c83 110 Vss 0.00128551f
c84 104 Vss 0.00368719f
c85 95 Vss 8.30816e-19
c86 94 Vss 0.00157211f
c87 93 Vss 8.30816e-19
c88 92 Vss 0.00157211f
c89 91 Vss 0.00860014f
c90 78 Vss 0.00407667f
c91 73 Vss 0.00419321f
c92 70 Vss 0.00352694f
c93 67 Vss 0.00278012f
c94 62 Vss 0.00185852f
c95 57 Vss 0.00149825f
c96 52 Vss 0.00105861f
c97 49 Vss 0.00997263f
c98 45 Vss 0.00798745f
c99 32 Vss 0.0350852f
c100 31 Vss 0.0994129f
c101 28 Vss 0.0350852f
c102 27 Vss 0.0994129f
c103 7 Vss 0.377882f
c104 3 Vss 0.379585f
r105 110 117 0.326018
r106 106 115 0.494161
r107 105 114 0.494161
r108 104 117 0.326018
r109 104 105 7.46046
r110 100 115 0.128424
r111 96 114 0.128424
r112 94 115 0.494161
r113 94 95 4.37625
r114 92 114 0.494161
r115 92 93 4.37625
r116 91 95 0.652036
r117 90 93 0.652036
r118 90 91 25.1739
r119 70 106 8.04396
r120 67 70 6.75193
r121 62 110 6.16843
r122 57 78 1.16709
r123 57 100 2.16729
r124 52 73 1.16709
r125 52 96 2.16729
r126 49 67 1.16709
r127 45 62 1.16709
r128 34 78 0.0476429
r129 32 34 1.45875
r130 31 38 0.652036
r131 31 34 1.45875
r132 30 73 0.0476429
r133 28 30 1.45875
r134 27 35 0.652036
r135 27 30 1.45875
r136 24 32 0.652036
r137 21 28 0.652036
r138 12 49 0.123773
r139 10 45 0.123773
r140 7 38 5.1348
r141 7 24 5.1348
r142 3 35 5.1348
r143 3 21 5.1348
.ends

.subckt PM_G4_MAJ3_N3_A 2 4 6 8 11 15 32 53 57 62 67 69 72 74 76 79 81 87 89 97
+ 100 109 Vss
c72 109 Vss 0.00544007f
c73 100 Vss 0.00497933f
c74 97 Vss 1.8079e-19
c75 94 Vss 7.63366e-19
c76 89 Vss 8.03875e-19
c77 87 Vss 8.73696e-19
c78 83 Vss 0.0024194f
c79 81 Vss 0.00445355f
c80 79 Vss 6.95023e-19
c81 76 Vss 0.00110877f
c82 75 Vss 0.00146569f
c83 74 Vss 0.00592189f
c84 69 Vss 0.00755424f
c85 67 Vss 0.0082356f
c86 62 Vss 0.00963114f
c87 57 Vss 0.135088f
c88 53 Vss 0.127963f
c89 32 Vss 0.217507f
c90 29 Vss 0.180502f
c91 27 Vss 0.0247918f
c92 11 Vss 1.44228f
c93 4 Vss 0.193588f
r94 109 112 0.1
r95 97 109 1.16709
r96 92 100 1.16709
r97 89 92 1.08364
r98 85 87 3.501
r99 84 97 0.0685365
r100 83 85 0.652036
r101 83 84 1.70882
r102 82 94 0.494161
r103 81 97 0.0685365
r104 81 82 7.46046
r105 77 94 0.128424
r106 77 79 3.501
r107 75 94 0.494161
r108 75 76 1.83386
r109 73 76 0.652036
r110 73 74 10.6697
r111 70 89 0.0685365
r112 70 72 1.41707
r113 69 74 0.652036
r114 69 72 8.79418
r115 67 87 1.16709
r116 62 79 1.16709
r117 55 57 4.53833
r118 52 112 0.0238214
r119 52 53 2.26917
r120 49 52 2.26917
r121 44 57 0.00605528
r122 43 53 0.00605528
r123 40 55 0.00605528
r124 39 49 0.00605528
r125 35 100 0.0476429
r126 33 35 0.326018
r127 33 35 0.1167
r128 32 36 0.652036
r129 32 35 6.7686
r130 29 100 0.357321
r131 27 35 0.326018
r132 27 29 0.40845
r133 15 44 5.1348
r134 15 40 5.1348
r135 11 15 17.9718
r136 11 43 5.1348
r137 11 15 17.9718
r138 11 39 5.1348
r139 8 67 0.123773
r140 6 62 0.123773
r141 4 36 5.1348
r142 2 29 4.72635
.ends

.subckt PM_G4_MAJ3_N3_BI 2 4 6 8 21 29 32 37 42 52 57 66 72 73 81 Vss
c58 81 Vss 5.35611e-19
c59 73 Vss 2.99365e-19
c60 72 Vss 7.27663e-19
c61 66 Vss 0.00156866f
c62 57 Vss 0.00147096f
c63 52 Vss 0.00166247f
c64 42 Vss 0.00166542f
c65 37 Vss 0.005464f
c66 32 Vss 0.00219142f
c67 29 Vss 0.00514303f
c68 21 Vss 0.166484f
c69 6 Vss 0.166484f
c70 4 Vss 0.00143493f
r71 77 81 0.655813
r72 72 73 0.65228
r73 71 72 3.42052
r74 66 71 0.65409
r75 42 57 1.16709
r76 42 73 2.1395
r77 37 52 1.16709
r78 37 81 12.0712
r79 37 66 1.96931
r80 32 49 1.16709
r81 32 77 3.25093
r82 29 49 0.1
r83 21 57 0.50025
r84 18 52 0.50025
r85 8 21 4.37625
r86 6 18 4.37625
r87 4 29 0.123773
r88 2 29 0.123773
.ends

.subckt PM_G4_MAJ3_N3_AI 2 4 7 11 31 37 43 46 51 60 69 Vss
c43 69 Vss 4.20376e-19
c44 60 Vss 0.00685099f
c45 51 Vss 0.00640177f
c46 46 Vss 9.78141e-19
c47 43 Vss 0.00452529f
c48 37 Vss 0.12791f
c49 31 Vss 0.134433f
c50 7 Vss 1.43419f
c51 4 Vss 0.00143493f
r52 65 69 0.652036
r53 60 63 0.1
r54 51 63 1.16709
r55 51 69 13.7539
r56 46 65 3.501
r57 43 46 1.16709
r58 36 60 0.0238214
r59 36 37 2.334
r60 33 36 2.20433
r61 29 31 4.53833
r62 26 37 0.00605528
r63 25 31 0.00605528
r64 22 33 0.00605528
r65 21 29 0.00605528
r66 11 26 5.1348
r67 11 22 5.1348
r68 7 11 17.9718
r69 7 25 5.1348
r70 7 11 17.9718
r71 7 21 5.1348
r72 4 43 0.123773
r73 2 43 0.123773
.ends

.subckt PM_G4_MAJ3_N3_B 2 4 6 8 16 17 26 38 42 45 50 55 60 65 73 74 80 87 92 93
+ Vss
c63 93 Vss 4.8362e-19
c64 92 Vss 0.00212566f
c65 87 Vss 9.92513e-19
c66 80 Vss 6.85439e-19
c67 74 Vss 5.17886e-19
c68 73 Vss 0.00375307f
c69 65 Vss 0.00163151f
c70 60 Vss 0.00118605f
c71 55 Vss 0.00132948f
c72 50 Vss 0.00183658f
c73 45 Vss 7.01705e-19
c74 38 Vss 0.00124968f
c75 26 Vss 0.166484f
c76 20 Vss 0.0247918f
c77 17 Vss 0.0349747f
c78 16 Vss 0.185505f
c79 8 Vss 0.166484f
c80 4 Vss 0.180512f
c81 2 Vss 0.192541f
r82 91 93 0.65409
r83 91 92 3.42052
r84 87 92 0.65228
r85 83 87 2.1006
r86 80 83 2.04225
r87 73 80 0.0685365
r88 73 74 10.3363
r89 69 74 0.652036
r90 50 65 1.16709
r91 50 93 2.00578
r92 45 60 1.16709
r93 45 83 0.0416786
r94 38 55 1.16709
r95 38 69 1.66714
r96 38 42 0.0833571
r97 36 55 0.238214
r98 33 65 0.50025
r99 26 60 0.50025
r100 24 36 0.262036
r101 20 36 0.326018
r102 20 24 0.05835
r103 17 36 6.7686
r104 16 36 0.326018
r105 16 36 0.1167
r106 13 17 0.652036
r107 8 33 4.37625
r108 6 26 4.37625
r109 4 24 5.07645
r110 2 13 5.1348
.ends

.subckt PM_G4_MAJ3_N3_C 2 4 12 17 20 25 51 Vss
c18 25 Vss 0.0055264f
c19 20 Vss 6.62222e-19
c20 17 Vss 0.00968607f
c21 12 Vss 0.00811861f
r22 25 51 1.89637
r23 20 51 8.169
r24 17 25 1.16709
r25 12 20 1.16709
r26 4 17 0.123773
r27 2 12 0.123773
.ends

.subckt PM_G4_MAJ3_N3_Z 2 4 6 8 23 27 30 33 Vss
c31 30 Vss 0.00306612f
c32 27 Vss 0.00807893f
c33 23 Vss 0.00720868f
c34 8 Vss 0.00143493f
c35 6 Vss 0.00143493f
r36 33 35 11.4616
r37 30 33 1.37539
r38 27 35 1.16709
r39 23 30 1.16709
r40 8 27 0.123773
r41 6 23 0.123773
r42 4 27 0.123773
r43 2 23 0.123773
.ends

.subckt G4_MAJ3_N3  VDD VSS A B C Z
*
* Z	Z
* C	C
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI19.X0 N_BI_XI19.X0_D N_VSS_XI19.X0_PGD N_B_XI19.X0_CG N_VSS_XI19.X0_PGD
+ N_VDD_XI19.X0_S TIGFET_HPNW12
XI18.X0 N_AI_XI18.X0_D N_VSS_XI18.X0_PGD N_A_XI18.X0_CG N_VSS_XI18.X0_PGD
+ N_VDD_XI18.X0_S TIGFET_HPNW12
XI17.X0 N_BI_XI17.X0_D N_VDD_XI17.X0_PGD N_B_XI17.X0_CG N_VDD_XI17.X0_PGD
+ N_VSS_XI17.X0_S TIGFET_HPNW12
XI16.X0 N_AI_XI16.X0_D N_VDD_XI16.X0_PGD N_A_XI16.X0_CG N_VDD_XI16.X0_PGD
+ N_VSS_XI16.X0_S TIGFET_HPNW12
XI22.X0 N_Z_XI22.X0_D N_AI_XI22.X0_PGD N_BI_XI22.X0_CG N_AI_XI22.X0_PGD
+ N_A_XI22.X0_S TIGFET_HPNW12
XI21.X0 N_Z_XI21.X0_D N_AI_XI21.X0_PGD N_B_XI21.X0_CG N_AI_XI21.X0_PGD
+ N_C_XI21.X0_S TIGFET_HPNW12
XI23.X0 N_Z_XI23.X0_D N_A_XI23.X0_PGD N_B_XI23.X0_CG N_A_XI23.X0_PGD
+ N_A_XI23.X0_S TIGFET_HPNW12
XI20.X0 N_Z_XI20.X0_D N_A_XI20.X0_PGD N_BI_XI20.X0_CG N_A_XI20.X0_PGD
+ N_C_XI20.X0_S TIGFET_HPNW12
*
x_PM_G4_MAJ3_N3_VDD N_VDD_XI19.X0_S N_VDD_XI18.X0_S N_VDD_XI17.X0_PGD
+ N_VDD_XI16.X0_PGD N_VDD_c_62_p N_VDD_c_4_p N_VDD_c_74_p N_VDD_c_63_p
+ N_VDD_c_8_p N_VDD_c_55_p N_VDD_c_64_p N_VDD_c_6_p N_VDD_c_33_p N_VDD_c_3_p
+ N_VDD_c_5_p N_VDD_c_39_p N_VDD_c_38_p VDD N_VDD_c_40_p N_VDD_c_9_p
+ N_VDD_c_42_p N_VDD_c_13_p N_VDD_c_17_p N_VDD_c_35_p N_VDD_c_36_p N_VDD_c_14_p
+ N_VDD_c_18_p Vss PM_G4_MAJ3_N3_VDD
x_PM_G4_MAJ3_N3_VSS N_VSS_XI19.X0_PGD N_VSS_XI18.X0_PGD N_VSS_XI17.X0_S
+ N_VSS_XI16.X0_S N_VSS_c_80_n N_VSS_c_82_n N_VSS_c_84_n N_VSS_c_86_n
+ N_VSS_c_123_p N_VSS_c_125_p N_VSS_c_87_n N_VSS_c_91_n N_VSS_c_95_n
+ N_VSS_c_96_n N_VSS_c_99_n N_VSS_c_100_n N_VSS_c_104_n N_VSS_c_108_n
+ N_VSS_c_113_n N_VSS_c_115_n N_VSS_c_116_n N_VSS_c_118_n N_VSS_c_119_n
+ N_VSS_c_120_n N_VSS_c_121_n VSS Vss PM_G4_MAJ3_N3_VSS
x_PM_G4_MAJ3_N3_A N_A_XI18.X0_CG N_A_XI16.X0_CG N_A_XI22.X0_S N_A_XI23.X0_S
+ N_A_XI23.X0_PGD N_A_XI20.X0_PGD N_A_c_158_n N_A_c_193_p N_A_c_195_p
+ N_A_c_168_n N_A_c_219_p N_A_c_159_n A N_A_c_174_n N_A_c_163_n N_A_c_214_p
+ N_A_c_180_p N_A_c_222_p N_A_c_165_n N_A_c_206_p N_A_c_166_n N_A_c_207_p Vss
+ PM_G4_MAJ3_N3_A
x_PM_G4_MAJ3_N3_BI N_BI_XI19.X0_D N_BI_XI17.X0_D N_BI_XI22.X0_CG N_BI_XI20.X0_CG
+ N_BI_c_243_n N_BI_c_230_n N_BI_c_232_n N_BI_c_240_n N_BI_c_260_p N_BI_c_248_n
+ N_BI_c_249_n N_BI_c_250_n N_BI_c_271_p N_BI_c_274_p N_BI_c_251_n Vss
+ PM_G4_MAJ3_N3_BI
x_PM_G4_MAJ3_N3_AI N_AI_XI18.X0_D N_AI_XI16.X0_D N_AI_XI22.X0_PGD
+ N_AI_XI21.X0_PGD N_AI_c_290_n N_AI_c_291_n N_AI_c_292_n N_AI_c_295_n
+ N_AI_c_299_n N_AI_c_308_n N_AI_c_309_n Vss PM_G4_MAJ3_N3_AI
x_PM_G4_MAJ3_N3_B N_B_XI19.X0_CG N_B_XI17.X0_CG N_B_XI21.X0_CG N_B_XI23.X0_CG
+ N_B_c_332_n N_B_c_342_n N_B_c_380_n N_B_c_333_n B N_B_c_360_n N_B_c_345_n
+ N_B_c_348_n N_B_c_365_n N_B_c_350_n N_B_c_338_n N_B_c_356_n N_B_c_357_n
+ N_B_c_374_n N_B_c_377_n N_B_c_378_n Vss PM_G4_MAJ3_N3_B
x_PM_G4_MAJ3_N3_C N_C_XI21.X0_S N_C_XI20.X0_S N_C_c_394_n N_C_c_407_p
+ N_C_c_395_n N_C_c_397_n C Vss PM_G4_MAJ3_N3_C
x_PM_G4_MAJ3_N3_Z N_Z_XI22.X0_D N_Z_XI21.X0_D N_Z_XI23.X0_D N_Z_XI20.X0_D
+ N_Z_c_412_n N_Z_c_437_n N_Z_c_417_n Z Vss PM_G4_MAJ3_N3_Z
cc_1 N_VDD_XI17.X0_PGD N_VSS_XI19.X0_PGD 0.00200629f
cc_2 N_VDD_XI16.X0_PGD N_VSS_XI18.X0_PGD 0.00200315f
cc_3 N_VDD_c_3_p N_VSS_XI18.X0_PGD 3.80615e-19
cc_4 N_VDD_c_4_p N_VSS_c_80_n 0.00200629f
cc_5 N_VDD_c_5_p N_VSS_c_80_n 3.89167e-19
cc_6 N_VDD_c_6_p N_VSS_c_82_n 3.80615e-19
cc_7 N_VDD_c_5_p N_VSS_c_82_n 3.89167e-19
cc_8 N_VDD_c_8_p N_VSS_c_84_n 0.00200315f
cc_9 N_VDD_c_9_p N_VSS_c_84_n 3.00203e-19
cc_10 N_VDD_c_9_p N_VSS_c_86_n 3.89167e-19
cc_11 N_VDD_c_6_p N_VSS_c_87_n 4.35319e-19
cc_12 N_VDD_c_5_p N_VSS_c_87_n 0.00141228f
cc_13 N_VDD_c_13_p N_VSS_c_87_n 9.22325e-19
cc_14 N_VDD_c_14_p N_VSS_c_87_n 3.48267e-19
cc_15 N_VDD_c_3_p N_VSS_c_91_n 4.35319e-19
cc_16 N_VDD_c_9_p N_VSS_c_91_n 0.00141228f
cc_17 N_VDD_c_17_p N_VSS_c_91_n 8.59637e-19
cc_18 N_VDD_c_18_p N_VSS_c_91_n 3.48267e-19
cc_19 N_VDD_c_13_p N_VSS_c_95_n 8.49247e-19
cc_20 N_VDD_XI16.X0_PGD N_VSS_c_96_n 2.8629e-19
cc_21 N_VDD_c_17_p N_VSS_c_96_n 0.00515616f
cc_22 N_VDD_c_18_p N_VSS_c_96_n 9.58524e-19
cc_23 N_VDD_c_9_p N_VSS_c_99_n 0.00403878f
cc_24 N_VDD_c_6_p N_VSS_c_100_n 3.66936e-19
cc_25 N_VDD_c_5_p N_VSS_c_100_n 0.00114511f
cc_26 N_VDD_c_13_p N_VSS_c_100_n 3.99794e-19
cc_27 N_VDD_c_14_p N_VSS_c_100_n 6.489e-19
cc_28 N_VDD_c_3_p N_VSS_c_104_n 3.66936e-19
cc_29 N_VDD_c_9_p N_VSS_c_104_n 0.00114511f
cc_30 N_VDD_c_17_p N_VSS_c_104_n 3.99794e-19
cc_31 N_VDD_c_18_p N_VSS_c_104_n 6.489e-19
cc_32 N_VDD_c_6_p N_VSS_c_108_n 0.00412661f
cc_33 N_VDD_c_33_p N_VSS_c_108_n 0.00936637f
cc_34 N_VDD_c_3_p N_VSS_c_108_n 0.00380969f
cc_35 N_VDD_c_35_p N_VSS_c_108_n 0.00104624f
cc_36 N_VDD_c_36_p N_VSS_c_108_n 0.0010706f
cc_37 N_VDD_c_5_p N_VSS_c_113_n 0.00331675f
cc_38 N_VDD_c_38_p N_VSS_c_113_n 2.97469e-19
cc_39 N_VDD_c_39_p N_VSS_c_115_n 0.00106807f
cc_40 N_VDD_c_40_p N_VSS_c_116_n 2.97469e-19
cc_41 N_VDD_c_9_p N_VSS_c_116_n 0.00331675f
cc_42 N_VDD_c_42_p N_VSS_c_118_n 0.00106807f
cc_43 N_VDD_c_5_p N_VSS_c_119_n 0.00602033f
cc_44 N_VDD_c_5_p N_VSS_c_120_n 7.74609e-19
cc_45 N_VDD_c_9_p N_VSS_c_121_n 7.74609e-19
cc_46 N_VDD_XI16.X0_PGD N_A_c_158_n 3.96972e-19
cc_47 N_VDD_XI16.X0_PGD N_A_c_159_n 5.06189e-19
cc_48 N_VDD_c_9_p N_A_c_159_n 2.07512e-19
cc_49 N_VDD_c_17_p N_A_c_159_n 2.39252e-19
cc_50 N_VDD_c_18_p N_A_c_159_n 2.01254e-19
cc_51 N_VDD_c_13_p N_A_c_163_n 5.45323e-19
cc_52 N_VDD_c_14_p N_A_c_163_n 4.10732e-19
cc_53 N_VDD_c_33_p N_A_c_165_n 9.17955e-19
cc_54 N_VDD_c_33_p N_A_c_166_n 5.22471e-19
cc_55 N_VDD_c_55_p N_BI_c_230_n 3.43419e-19
cc_56 N_VDD_c_38_p N_BI_c_230_n 3.72199e-19
cc_57 N_VDD_c_55_p N_BI_c_232_n 3.48267e-19
cc_58 N_VDD_c_5_p N_BI_c_232_n 3.12875e-19
cc_59 N_VDD_c_38_p N_BI_c_232_n 5.2846e-19
cc_60 N_VDD_XI17.X0_PGD N_AI_XI22.X0_PGD 2.84861e-19
cc_61 N_VDD_XI16.X0_PGD N_AI_XI22.X0_PGD 3.10667e-19
cc_62 N_VDD_c_62_p N_AI_c_290_n 2.84861e-19
cc_63 N_VDD_c_63_p N_AI_c_291_n 3.10667e-19
cc_64 N_VDD_c_64_p N_AI_c_292_n 3.43419e-19
cc_65 N_VDD_c_40_p N_AI_c_292_n 3.72199e-19
cc_66 N_VDD_c_9_p N_AI_c_292_n 2.74986e-19
cc_67 N_VDD_c_64_p N_AI_c_295_n 3.48267e-19
cc_68 N_VDD_c_3_p N_AI_c_295_n 2.34601e-19
cc_69 N_VDD_c_40_p N_AI_c_295_n 5.226e-19
cc_70 N_VDD_c_9_p N_AI_c_295_n 2.9533e-19
cc_71 N_VDD_c_17_p N_AI_c_299_n 9.90259e-19
cc_72 N_VDD_c_33_p N_B_XI19.X0_CG 3.68219e-19
cc_73 N_VDD_XI17.X0_PGD N_B_c_332_n 4.01605e-19
cc_74 N_VDD_c_74_p N_B_c_333_n 2.01616e-19
cc_75 N_VDD_c_33_p N_B_c_333_n 3.58277e-19
cc_76 N_VDD_c_14_p N_B_c_333_n 2.07877e-19
cc_77 N_VSS_XI18.X0_PGD N_A_c_158_n 3.96972e-19
cc_78 N_VSS_c_123_p N_A_c_168_n 3.43419e-19
cc_79 N_VSS_c_123_p N_A_c_159_n 2.21087e-19
cc_80 N_VSS_c_125_p N_A_c_159_n 4.13509e-19
cc_81 N_VSS_c_95_n N_A_c_159_n 2.50981e-19
cc_82 N_VSS_c_96_n N_A_c_159_n 7.05313e-19
cc_83 N_VSS_c_99_n N_A_c_159_n 2.62883e-19
cc_84 N_VSS_c_123_p N_A_c_174_n 9.18655e-19
cc_85 N_VSS_c_95_n N_A_c_174_n 0.00202874f
cc_86 N_VSS_c_95_n N_A_c_163_n 0.00196507f
cc_87 N_VSS_c_104_n N_A_c_165_n 4.60155e-19
cc_88 N_VSS_c_108_n N_A_c_165_n 5.04162e-19
cc_89 N_VSS_c_91_n N_A_c_166_n 2.15082e-19
cc_90 N_VSS_c_123_p N_BI_c_230_n 3.43419e-19
cc_91 N_VSS_c_123_p N_BI_c_232_n 3.48267e-19
cc_92 N_VSS_c_95_n N_BI_c_232_n 0.00105024f
cc_93 N_VSS_c_108_n N_BI_c_232_n 0.00120568f
cc_94 N_VSS_c_119_n N_BI_c_232_n 2.38659e-19
cc_95 N_VSS_c_95_n N_BI_c_240_n 4.33962e-19
cc_96 N_VSS_c_119_n N_BI_c_240_n 6.35155e-19
cc_97 N_VSS_c_125_p N_AI_c_292_n 3.43419e-19
cc_98 N_VSS_c_96_n N_AI_c_292_n 3.48267e-19
cc_99 N_VSS_c_125_p N_AI_c_295_n 3.48267e-19
cc_100 N_VSS_c_91_n N_AI_c_295_n 0.00173332f
cc_101 N_VSS_c_96_n N_AI_c_295_n 0.00178201f
cc_102 N_VSS_c_108_n N_AI_c_295_n 0.00136931f
cc_103 N_VSS_c_96_n N_AI_c_299_n 0.00200998f
cc_104 N_VSS_c_99_n N_AI_c_299_n 0.00674978f
cc_105 N_VSS_c_96_n N_AI_c_308_n 2.82216e-19
cc_106 N_VSS_c_99_n N_AI_c_309_n 0.00178766f
cc_107 N_VSS_XI19.X0_PGD N_B_c_332_n 4.01605e-19
cc_108 N_VSS_c_108_n N_B_c_333_n 7.40204e-19
cc_109 N_VSS_c_95_n N_B_c_338_n 4.25717e-19
cc_110 N_VSS_c_125_p N_C_c_394_n 3.43419e-19
cc_111 N_VSS_c_125_p N_C_c_395_n 3.48267e-19
cc_112 N_VSS_c_96_n N_C_c_395_n 6.01757e-19
cc_113 N_A_c_180_p N_BI_XI22.X0_CG 2.10479e-19
cc_114 N_A_XI23.X0_PGD N_BI_c_243_n 9.65637e-19
cc_115 N_A_c_159_n N_BI_c_232_n 3.45962e-19
cc_116 N_A_c_174_n N_BI_c_232_n 5.71688e-19
cc_117 N_A_c_174_n N_BI_c_240_n 0.00169296f
cc_118 N_A_c_180_p N_BI_c_240_n 6.66847e-19
cc_119 N_A_c_174_n N_BI_c_248_n 3.37713e-19
cc_120 N_A_XI23.X0_PGD N_BI_c_249_n 0.00245019f
cc_121 N_A_c_180_p N_BI_c_250_n 9.24697e-19
cc_122 N_A_c_159_n N_BI_c_251_n 8.09947e-19
cc_123 N_A_XI23.X0_PGD N_AI_XI22.X0_PGD 0.0174035f
cc_124 N_A_c_174_n N_AI_XI22.X0_PGD 8.23587e-19
cc_125 N_A_c_180_p N_AI_XI22.X0_PGD 9.89767e-19
cc_126 N_A_c_193_p N_AI_c_290_n 0.00196311f
cc_127 N_A_c_180_p N_AI_c_290_n 0.00103585f
cc_128 N_A_c_195_p N_AI_c_291_n 0.00200674f
cc_129 N_A_c_158_n N_AI_c_292_n 6.90199e-19
cc_130 N_A_c_159_n N_AI_c_295_n 5.79974e-19
cc_131 N_A_c_159_n N_AI_c_299_n 0.00132412f
cc_132 N_A_XI23.X0_PGD N_B_XI23.X0_CG 9.65637e-19
cc_133 N_A_c_158_n N_B_c_332_n 0.0036037f
cc_134 N_A_c_159_n N_B_c_332_n 8.51862e-19
cc_135 N_A_c_166_n N_B_c_342_n 6.91203e-19
cc_136 N_A_c_159_n N_B_c_333_n 0.00120731f
cc_137 N_A_c_174_n N_B_c_333_n 0.00118668f
cc_138 N_A_c_180_p N_B_c_345_n 3.57869e-19
cc_139 N_A_c_206_p N_B_c_345_n 3.46877e-19
cc_140 N_A_c_207_p N_B_c_345_n 2.26741e-19
cc_141 N_A_c_159_n N_B_c_348_n 7.40468e-19
cc_142 N_A_c_174_n N_B_c_348_n 5.93411e-19
cc_143 N_A_XI23.X0_PGD N_B_c_350_n 0.00312702f
cc_144 N_A_c_206_p N_B_c_350_n 2.30774e-19
cc_145 N_A_c_159_n N_B_c_338_n 0.00230073f
cc_146 N_A_c_174_n N_B_c_338_n 0.00203212f
cc_147 N_A_c_214_p N_B_c_338_n 3.55185e-19
cc_148 N_A_c_180_p N_B_c_338_n 4.84888e-19
cc_149 N_A_c_159_n N_B_c_356_n 4.20277e-19
cc_150 N_A_c_159_n N_B_c_357_n 2.29222e-19
cc_151 N_A_c_168_n N_Z_c_412_n 3.43419e-19
cc_152 N_A_c_219_p N_Z_c_412_n 3.43419e-19
cc_153 N_A_c_214_p N_Z_c_412_n 3.48267e-19
cc_154 N_A_c_180_p N_Z_c_412_n 5.52794e-19
cc_155 N_A_c_222_p N_Z_c_412_n 3.48267e-19
cc_156 N_A_XI23.X0_PGD N_Z_c_417_n 6.68421e-19
cc_157 N_A_c_168_n N_Z_c_417_n 3.48267e-19
cc_158 N_A_c_219_p N_Z_c_417_n 3.48267e-19
cc_159 N_A_c_174_n N_Z_c_417_n 0.00158522f
cc_160 N_A_c_214_p N_Z_c_417_n 7.9714e-19
cc_161 N_A_c_180_p N_Z_c_417_n 9.31302e-19
cc_162 N_A_c_222_p N_Z_c_417_n 8.16241e-19
cc_163 N_BI_XI22.X0_CG N_AI_XI22.X0_PGD 9.47088e-19
cc_164 N_BI_c_248_n N_AI_XI22.X0_PGD 0.00312702f
cc_165 N_BI_c_251_n N_AI_c_295_n 2.92168e-19
cc_166 N_BI_c_240_n N_AI_c_299_n 3.11073e-19
cc_167 N_BI_c_230_n N_B_c_332_n 6.90199e-19
cc_168 N_BI_c_240_n N_B_c_333_n 0.0014575f
cc_169 N_BI_c_240_n N_B_c_360_n 6.83975e-19
cc_170 N_BI_c_248_n N_B_c_360_n 4.99367e-19
cc_171 N_BI_c_260_p N_B_c_345_n 0.0018485f
cc_172 N_BI_c_249_n N_B_c_345_n 4.99367e-19
cc_173 N_BI_c_250_n N_B_c_345_n 0.00165504f
cc_174 N_BI_c_248_n N_B_c_365_n 0.00521054f
cc_175 N_BI_c_249_n N_B_c_365_n 7.2092e-19
cc_176 N_BI_c_260_p N_B_c_350_n 4.99367e-19
cc_177 N_BI_c_248_n N_B_c_350_n 6.22265e-19
cc_178 N_BI_c_249_n N_B_c_350_n 0.00494884f
cc_179 N_BI_c_240_n N_B_c_338_n 0.00536154f
cc_180 N_BI_c_240_n N_B_c_357_n 2.67017e-19
cc_181 N_BI_c_250_n N_B_c_357_n 0.0013533f
cc_182 N_BI_c_271_p N_B_c_357_n 0.00340518f
cc_183 N_BI_c_240_n N_B_c_374_n 4.99817e-19
cc_184 N_BI_c_250_n N_B_c_374_n 9.84686e-19
cc_185 N_BI_c_274_p N_B_c_374_n 7.60478e-19
cc_186 N_BI_c_271_p N_B_c_377_n 0.00181541f
cc_187 N_BI_c_240_n N_B_c_378_n 0.00145553f
cc_188 N_BI_c_250_n N_B_c_378_n 8.77567e-19
cc_189 N_BI_c_240_n N_C_c_397_n 9.46412e-19
cc_190 N_BI_c_260_p N_C_c_397_n 0.00112215f
cc_191 N_BI_c_274_p N_C_c_397_n 2.41224e-19
cc_192 N_BI_c_240_n N_Z_c_417_n 0.00190811f
cc_193 N_BI_c_260_p N_Z_c_417_n 0.00192905f
cc_194 N_BI_c_248_n N_Z_c_417_n 8.66889e-19
cc_195 N_BI_c_249_n N_Z_c_417_n 8.66889e-19
cc_196 N_BI_c_250_n N_Z_c_417_n 0.00108781f
cc_197 N_BI_c_271_p N_Z_c_417_n 0.00210701f
cc_198 N_BI_c_274_p N_Z_c_417_n 0.00102097f
cc_199 N_AI_XI22.X0_PGD N_B_c_380_n 9.65637e-19
cc_200 N_AI_c_299_n N_B_c_360_n 3.12862e-19
cc_201 N_AI_c_308_n N_B_c_360_n 2.26741e-19
cc_202 N_AI_XI22.X0_PGD N_B_c_365_n 0.00312702f
cc_203 N_AI_c_299_n N_B_c_338_n 0.00252591f
cc_204 N_AI_c_299_n N_C_c_395_n 0.00111024f
cc_205 N_AI_c_299_n N_C_c_397_n 0.0016345f
cc_206 N_AI_XI22.X0_PGD N_Z_c_417_n 3.73496e-19
cc_207 N_B_c_338_n N_C_c_395_n 4.14759e-19
cc_208 N_B_c_345_n N_C_c_397_n 8.23684e-19
cc_209 N_B_c_338_n N_C_c_397_n 3.71981e-19
cc_210 N_B_c_374_n N_C_c_397_n 0.0032187f
cc_211 N_B_c_360_n N_Z_c_417_n 0.00192136f
cc_212 N_B_c_345_n N_Z_c_417_n 0.0019232f
cc_213 N_B_c_365_n N_Z_c_417_n 8.66889e-19
cc_214 N_B_c_350_n N_Z_c_417_n 8.66889e-19
cc_215 N_B_c_357_n N_Z_c_417_n 4.75654e-19
cc_216 N_C_c_394_n N_Z_c_437_n 3.43419e-19
cc_217 N_C_c_407_p N_Z_c_437_n 3.43419e-19
cc_218 N_C_c_395_n N_Z_c_437_n 3.48267e-19
cc_219 N_C_c_397_n N_Z_c_437_n 3.48267e-19
cc_220 N_C_c_395_n N_Z_c_417_n 6.20216e-19
cc_221 N_C_c_397_n N_Z_c_417_n 0.00134739f
*
.ends
*
*
.subckt MAJ3_HPNW12 A B C Y VDD VSS
xgate (VDD VSS A B C Y) G4_MAJ3_N3
.ends
*
* File: G3_MIN3_T6_N3.pex.netlist
* Created: Mon Apr  4 15:49:45 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MIN3_T6_N3_VSS 2 4 6 8 10 12 27 32 37 40 42 45 53 57 60 65 70 75
+ 88 89 93 99 101 106 109 Vss
c64 107 Vss 6.47574e-19
c65 106 Vss 0.00464148f
c66 101 Vss 0.00213175f
c67 99 Vss 0.0082833f
c68 94 Vss 0.00138375f
c69 93 Vss 0.00819383f
c70 89 Vss 6.61473e-19
c71 88 Vss 0.0060976f
c72 75 Vss 0.006288f
c73 70 Vss 1.73335e-19
c74 65 Vss 0.00209248f
c75 60 Vss 0.00138481f
c76 57 Vss 0.0103194f
c77 53 Vss 0.00454903f
c78 45 Vss 0.0856842f
c79 42 Vss 0.0855647f
c80 37 Vss 0.0648277f
c81 32 Vss 0.103906f
c82 27 Vss 0.306999f
c83 22 Vss 0.141041f
c84 10 Vss 0.186558f
c85 8 Vss 0.00171982f
c86 6 Vss 0.188337f
c87 2 Vss 0.185627f
r88 106 109 0.326018
r89 105 106 5.50157
r90 101 105 0.655813
r91 100 107 0.494161
r92 99 109 0.326018
r93 99 100 13.0037
r94 95 107 0.128424
r95 93 107 0.494161
r96 93 94 10.0862
r97 88 94 0.652036
r98 87 89 0.655813
r99 87 88 16.4214
r100 70 101 1.82344
r101 65 95 6.16843
r102 60 75 1.16709
r103 60 89 1.82344
r104 57 70 1.16709
r105 53 65 1.16709
r106 45 47 1.8672
r107 42 44 1.8672
r108 40 75 0.50025
r109 37 40 1.92555
r110 33 47 0.0685365
r111 32 34 0.652036
r112 32 33 2.8008
r113 29 47 0.5835
r114 28 42 0.0685365
r115 27 45 0.0685365
r116 27 28 10.9698
r117 24 44 0.5835
r118 23 37 0.0685365
r119 22 44 0.0685365
r120 22 23 4.7847
r121 12 57 0.123773
r122 10 34 5.1348
r123 8 53 0.123773
r124 6 29 5.1348
r125 4 53 0.123773
r126 2 24 5.1348
.ends

.subckt PM_G3_MIN3_T6_N3_VDD 2 4 6 8 10 12 27 32 42 45 53 57 60 61 63 65 69 71
+ 73 78 81 83 Vss
c74 83 Vss 0.00747336f
c75 79 Vss 7.84502e-19
c76 78 Vss 0.00603664f
c77 73 Vss 0.00149586f
c78 71 Vss 0.0125181f
c79 69 Vss 0.00223179f
c80 65 Vss 0.00180228f
c81 63 Vss 7.51405e-19
c82 62 Vss 0.00180268f
c83 61 Vss 0.00800879f
c84 60 Vss 0.00954496f
c85 57 Vss 0.00979559f
c86 53 Vss 0.00450493f
c87 45 Vss 0.0849231f
c88 42 Vss 0.0854945f
c89 38 Vss 0.0711342f
c90 32 Vss 0.106731f
c91 27 Vss 0.308123f
c92 22 Vss 0.144485f
c93 12 Vss 0.187032f
c94 8 Vss 0.187847f
c95 6 Vss 0.00171982f
c96 4 Vss 0.18764f
r97 78 81 0.349767
r98 77 78 5.50157
r99 73 81 0.306046
r100 73 75 1.82344
r101 72 79 0.494161
r102 71 77 0.652036
r103 71 72 13.0037
r104 67 79 0.128424
r105 67 69 6.16843
r106 65 83 1.16709
r107 63 65 1.82344
r108 61 79 0.494161
r109 61 62 10.0862
r110 60 63 0.655813
r111 59 62 0.652036
r112 59 60 16.4214
r113 57 75 1.16709
r114 53 69 1.16709
r115 45 46 1.8672
r116 42 43 1.8672
r117 38 83 0.50025
r118 38 40 1.92555
r119 33 45 0.0685365
r120 32 34 0.652036
r121 32 33 2.8008
r122 29 45 0.5835
r123 28 43 0.0685365
r124 27 46 0.0685365
r125 27 28 10.9698
r126 24 42 0.5835
r127 23 40 0.0685365
r128 22 42 0.0685365
r129 22 23 4.7847
r130 12 34 5.1348
r131 10 57 0.123773
r132 8 29 5.1348
r133 6 53 0.123773
r134 4 24 5.1348
r135 2 53 0.123773
.ends

.subckt PM_G3_MIN3_T6_N3_Z 2 4 6 8 10 12 32 36 41 45 49 53 55 59 63 67 Vss
c55 67 Vss 3.51451e-19
c56 65 Vss 2.45386e-19
c57 63 Vss 0.00102688f
c58 59 Vss 7.58182e-19
c59 55 Vss 0.0050105f
c60 53 Vss 6.51205e-19
c61 49 Vss 5.16244e-19
c62 45 Vss 0.00816234f
c63 41 Vss 0.00751221f
c64 36 Vss 0.00857712f
c65 32 Vss 0.00789336f
c66 12 Vss 0.00171982f
c67 10 Vss 0.00171982f
r68 61 67 0.494161
r69 61 63 3.95946
r70 57 67 0.494161
r71 57 59 3.95946
r72 56 65 0.128424
r73 55 67 0.128424
r74 55 56 10.3363
r75 51 65 0.494161
r76 51 53 3.95946
r77 47 65 0.494161
r78 47 49 3.95946
r79 45 63 1.16709
r80 41 59 1.16709
r81 36 53 1.16709
r82 32 49 1.16709
r83 12 45 0.123773
r84 10 41 0.123773
r85 8 45 0.123773
r86 6 41 0.123773
r87 4 36 0.123773
r88 2 32 0.123773
.ends

.subckt PM_G3_MIN3_T6_N3_C 2 4 6 8 14 20 26 33 38 43 Vss
c33 43 Vss 0.00462472f
c34 38 Vss 0.00103857f
c35 33 Vss 0.00642701f
c36 26 Vss 7.12876e-22
c37 20 Vss 0.486644f
c38 14 Vss 0.489687f
r39 33 43 1.16709
r40 29 38 1.16709
r41 29 33 11.5033
r42 26 29 0.166714
r43 20 43 0.50025
r44 14 38 0.50025
r45 6 8 12.7203
r46 6 20 4.37625
r47 2 4 12.7203
r48 2 14 4.37625
.ends

.subckt PM_G3_MIN3_T6_N3_B 2 4 6 8 17 18 26 29 32 35 Vss
c31 35 Vss 0.00167659f
c32 26 Vss 0.0837857f
c33 18 Vss 0.034641f
c34 17 Vss 0.09638f
c35 6 Vss 0.506992f
c36 2 Vss 0.554218f
r37 32 35 1.16709
r38 29 32 0.0729375
r39 24 35 0.0476429
r40 24 26 1.92555
r41 17 19 0.652036
r42 17 18 2.8008
r43 14 26 0.0685365
r44 13 18 0.652036
r45 6 8 12.7203
r46 6 19 5.1348
r47 4 14 5.1348
r48 2 4 12.7203
r49 2 13 5.1348
.ends

.subckt PM_G3_MIN3_T6_N3_A 2 4 6 8 17 29 34 38 41 46 Vss
c29 46 Vss 0.00528506f
c30 41 Vss 0.00159958f
c31 38 Vss 3.66482e-19
c32 34 Vss 0.00172621f
c33 29 Vss 3.54075e-22
c34 26 Vss 0.0871371f
c35 6 Vss 0.515115f
c36 2 Vss 0.485149f
r37 34 46 1.16709
r38 34 38 0.109406
r39 29 41 1.16709
r40 29 34 5.03269
r41 24 46 0.0476429
r42 24 26 1.92555
r43 19 26 0.0685365
r44 17 41 0.50025
r45 8 19 5.1348
r46 6 8 12.7203
r47 4 17 4.37625
r48 2 4 12.7203
.ends

.subckt G3_MIN3_T6_N3  VSS VDD Z C B A
*
* A	A
* B	B
* C	C
* Z	Z
* VDD	VDD
* VSS	VSS
XI24.X0 N_Z_XI24.X0_D N_VSS_XI24.X0_PGD N_C_XI24.X0_CG N_B_XI24.X0_PGS
+ N_VDD_XI24.X0_S TIGFET_HPNW12
XI20.X0 N_Z_XI20.X0_D N_VDD_XI20.X0_PGD N_C_XI20.X0_CG N_B_XI20.X0_PGS
+ N_VSS_XI20.X0_S TIGFET_HPNW12
XI23.X0 N_Z_XI23.X0_D N_VSS_XI23.X0_PGD N_A_XI23.X0_CG N_B_XI23.X0_PGS
+ N_VDD_XI23.X0_S TIGFET_HPNW12
XI22.X0 N_Z_XI22.X0_D N_VDD_XI22.X0_PGD N_A_XI22.X0_CG N_B_XI22.X0_PGS
+ N_VSS_XI22.X0_S TIGFET_HPNW12
XI25.X0 N_Z_XI25.X0_D N_VSS_XI25.X0_PGD N_C_XI25.X0_CG N_A_XI25.X0_PGS
+ N_VDD_XI25.X0_S TIGFET_HPNW12
XI21.X0 N_Z_XI21.X0_D N_VDD_XI21.X0_PGD N_C_XI21.X0_CG N_A_XI21.X0_PGS
+ N_VSS_XI21.X0_S TIGFET_HPNW12
*
x_PM_G3_MIN3_T6_N3_VSS N_VSS_XI24.X0_PGD N_VSS_XI20.X0_S N_VSS_XI23.X0_PGD
+ N_VSS_XI22.X0_S N_VSS_XI25.X0_PGD N_VSS_XI21.X0_S N_VSS_c_19_p N_VSS_c_22_p
+ N_VSS_c_6_p N_VSS_c_12_p N_VSS_c_13_p N_VSS_c_46_p N_VSS_c_4_p N_VSS_c_29_p
+ N_VSS_c_7_p N_VSS_c_17_p N_VSS_c_23_p N_VSS_c_8_p N_VSS_c_9_p N_VSS_c_10_p
+ N_VSS_c_18_p N_VSS_c_43_p N_VSS_c_24_p N_VSS_c_62_p VSS Vss
+ PM_G3_MIN3_T6_N3_VSS
x_PM_G3_MIN3_T6_N3_VDD N_VDD_XI24.X0_S N_VDD_XI20.X0_PGD N_VDD_XI23.X0_S
+ N_VDD_XI22.X0_PGD N_VDD_XI25.X0_S N_VDD_XI21.X0_PGD N_VDD_c_68_n N_VDD_c_137_p
+ N_VDD_c_130_p N_VDD_c_129_p N_VDD_c_69_n N_VDD_c_96_p N_VDD_c_70_n
+ N_VDD_c_75_n N_VDD_c_79_n N_VDD_c_80_n N_VDD_c_83_n N_VDD_c_85_n N_VDD_c_87_n
+ N_VDD_c_119_p VDD N_VDD_c_89_n Vss PM_G3_MIN3_T6_N3_VDD
x_PM_G3_MIN3_T6_N3_Z N_Z_XI24.X0_D N_Z_XI20.X0_D N_Z_XI23.X0_D N_Z_XI22.X0_D
+ N_Z_XI25.X0_D N_Z_XI21.X0_D N_Z_c_154_n N_Z_c_139_n N_Z_c_159_n N_Z_c_141_n
+ N_Z_c_145_n N_Z_c_146_n N_Z_c_149_n N_Z_c_172_n N_Z_c_151_n Z Vss
+ PM_G3_MIN3_T6_N3_Z
x_PM_G3_MIN3_T6_N3_C N_C_XI24.X0_CG N_C_XI20.X0_CG N_C_XI25.X0_CG N_C_XI21.X0_CG
+ N_C_c_194_n N_C_c_195_n C N_C_c_196_n N_C_c_197_n N_C_c_198_n Vss
+ PM_G3_MIN3_T6_N3_C
x_PM_G3_MIN3_T6_N3_B N_B_XI24.X0_PGS N_B_XI20.X0_PGS N_B_XI23.X0_PGS
+ N_B_XI22.X0_PGS N_B_c_231_n N_B_c_232_n N_B_c_240_n B N_B_c_234_n N_B_c_242_n
+ Vss PM_G3_MIN3_T6_N3_B
x_PM_G3_MIN3_T6_N3_A N_A_XI23.X0_CG N_A_XI22.X0_CG N_A_XI25.X0_PGS
+ N_A_XI21.X0_PGS N_A_c_274_n N_A_c_259_n N_A_c_261_n A N_A_c_269_n N_A_c_270_n
+ Vss PM_G3_MIN3_T6_N3_A
cc_1 N_VSS_XI24.X0_PGD N_VDD_XI20.X0_PGD 6.54383e-19
cc_2 N_VSS_XI23.X0_PGD N_VDD_XI22.X0_PGD 6.54383e-19
cc_3 N_VSS_XI25.X0_PGD N_VDD_XI21.X0_PGD 6.43556e-19
cc_4 N_VSS_c_4_p N_VDD_c_68_n 5.08814e-19
cc_5 N_VSS_c_4_p N_VDD_c_69_n 7.73686e-19
cc_6 N_VSS_c_6_p N_VDD_c_70_n 2.63314e-19
cc_7 N_VSS_c_7_p N_VDD_c_70_n 0.00161042f
cc_8 N_VSS_c_8_p N_VDD_c_70_n 0.00115993f
cc_9 N_VSS_c_9_p N_VDD_c_70_n 0.00777883f
cc_10 N_VSS_c_10_p N_VDD_c_70_n 0.00186982f
cc_11 N_VSS_c_6_p N_VDD_c_75_n 8.77582e-19
cc_12 N_VSS_c_12_p N_VDD_c_75_n 3.72495e-19
cc_13 N_VSS_c_13_p N_VDD_c_75_n 7.64639e-19
cc_14 N_VSS_c_7_p N_VDD_c_75_n 9.97468e-19
cc_15 N_VSS_c_9_p N_VDD_c_79_n 0.00179061f
cc_16 N_VSS_c_7_p N_VDD_c_80_n 3.76254e-19
cc_17 N_VSS_c_17_p N_VDD_c_80_n 2.77394e-19
cc_18 N_VSS_c_18_p N_VDD_c_80_n 4.66156e-19
cc_19 N_VSS_c_19_p N_VDD_c_83_n 0.00120485f
cc_20 N_VSS_c_7_p N_VDD_c_83_n 4.38149e-19
cc_21 N_VSS_c_19_p N_VDD_c_85_n 8.70027e-19
cc_22 N_VSS_c_22_p N_VDD_c_85_n 8.24361e-19
cc_23 N_VSS_c_23_p N_VDD_c_87_n 2.543e-19
cc_24 N_VSS_c_24_p N_VDD_c_87_n 0.00120656f
cc_25 N_VSS_c_8_p N_VDD_c_89_n 2.36483e-19
cc_26 N_VSS_c_4_p N_Z_c_139_n 3.43419e-19
cc_27 N_VSS_c_17_p N_Z_c_139_n 3.48267e-19
cc_28 N_VSS_c_4_p N_Z_c_141_n 3.43419e-19
cc_29 N_VSS_c_29_p N_Z_c_141_n 3.43419e-19
cc_30 N_VSS_c_17_p N_Z_c_141_n 3.48267e-19
cc_31 N_VSS_c_23_p N_Z_c_141_n 3.48267e-19
cc_32 N_VSS_c_9_p N_Z_c_145_n 0.00213783f
cc_33 N_VSS_c_4_p N_Z_c_146_n 3.48267e-19
cc_34 N_VSS_c_17_p N_Z_c_146_n 5.02484e-19
cc_35 N_VSS_c_18_p N_Z_c_146_n 4.85461e-19
cc_36 N_VSS_c_4_p N_Z_c_149_n 4.81023e-19
cc_37 N_VSS_c_17_p N_Z_c_149_n 6.34336e-19
cc_38 N_VSS_c_29_p N_Z_c_151_n 3.48267e-19
cc_39 N_VSS_c_17_p N_Z_c_151_n 5.37696e-19
cc_40 N_VSS_c_23_p N_Z_c_151_n 5.71987e-19
cc_41 N_VSS_XI24.X0_PGD N_C_c_194_n 4.30517e-19
cc_42 N_VSS_XI25.X0_PGD N_C_c_195_n 4.94554e-19
cc_43 N_VSS_c_43_p N_C_c_196_n 5.18193e-19
cc_44 N_VSS_XI24.X0_PGD N_C_c_197_n 4.3583e-19
cc_45 N_VSS_XI25.X0_PGD N_C_c_198_n 3.76133e-19
cc_46 N_VSS_c_46_p N_C_c_198_n 2.17009e-19
cc_47 N_VSS_XI24.X0_PGD N_B_XI24.X0_PGS 0.00109504f
cc_48 N_VSS_XI23.X0_PGD N_B_XI24.X0_PGS 2.15671e-19
cc_49 N_VSS_XI23.X0_PGD N_B_XI23.X0_PGS 0.00177732f
cc_50 N_VSS_XI25.X0_PGD N_B_XI23.X0_PGS 2.22194e-19
cc_51 N_VSS_c_46_p N_B_c_231_n 0.00177732f
cc_52 N_VSS_c_19_p N_B_c_232_n 0.00722404f
cc_53 N_VSS_c_13_p N_B_c_232_n 0.00109504f
cc_54 N_VSS_c_17_p N_B_c_234_n 2.11465e-19
cc_55 N_VSS_c_9_p N_B_c_234_n 2.74582e-19
cc_56 N_VSS_c_18_p N_B_c_234_n 4.28832e-19
cc_57 N_VSS_c_19_p N_A_XI23.X0_CG 2.64949e-19
cc_58 N_VSS_c_17_p N_A_c_259_n 3.13396e-19
cc_59 N_VSS_c_43_p N_A_c_259_n 5.88825e-19
cc_60 N_VSS_c_17_p N_A_c_261_n 0.00159318f
cc_61 N_VSS_c_43_p N_A_c_261_n 0.00925582f
cc_62 N_VSS_c_62_p N_A_c_261_n 7.74234e-19
cc_63 N_VSS_c_43_p A 5.88825e-19
cc_64 N_VSS_c_62_p A 3.28646e-19
cc_65 N_VDD_c_69_n N_Z_c_154_n 3.43419e-19
cc_66 N_VDD_c_70_n N_Z_c_154_n 3.70842e-19
cc_67 N_VDD_c_75_n N_Z_c_154_n 2.74986e-19
cc_68 N_VDD_c_83_n N_Z_c_154_n 3.48267e-19
cc_69 N_VDD_c_70_n N_Z_c_139_n 3.70842e-19
cc_70 N_VDD_c_69_n N_Z_c_159_n 3.43419e-19
cc_71 N_VDD_c_96_p N_Z_c_159_n 3.43419e-19
cc_72 N_VDD_c_83_n N_Z_c_159_n 3.48267e-19
cc_73 N_VDD_c_85_n N_Z_c_159_n 2.74986e-19
cc_74 N_VDD_c_87_n N_Z_c_159_n 3.72199e-19
cc_75 N_VDD_c_69_n N_Z_c_145_n 3.48267e-19
cc_76 N_VDD_c_70_n N_Z_c_145_n 0.00440367f
cc_77 N_VDD_c_75_n N_Z_c_145_n 5.29921e-19
cc_78 N_VDD_c_83_n N_Z_c_145_n 7.15874e-19
cc_79 N_VDD_c_69_n N_Z_c_149_n 4.81023e-19
cc_80 N_VDD_c_75_n N_Z_c_149_n 3.00455e-19
cc_81 N_VDD_c_83_n N_Z_c_149_n 8.48441e-19
cc_82 N_VDD_c_85_n N_Z_c_149_n 4.56827e-19
cc_83 N_VDD_c_69_n N_Z_c_172_n 3.48267e-19
cc_84 N_VDD_c_96_p N_Z_c_172_n 3.48267e-19
cc_85 N_VDD_c_83_n N_Z_c_172_n 7.23486e-19
cc_86 N_VDD_c_85_n N_Z_c_172_n 4.06373e-19
cc_87 N_VDD_c_87_n N_Z_c_172_n 8.5731e-19
cc_88 N_VDD_c_70_n C 2.30446e-19
cc_89 N_VDD_c_75_n C 0.00138543f
cc_90 N_VDD_c_83_n C 0.00115642f
cc_91 N_VDD_c_75_n N_C_c_196_n 7.64872e-19
cc_92 N_VDD_c_83_n N_C_c_196_n 0.00221688f
cc_93 N_VDD_c_85_n N_C_c_196_n 0.0053512f
cc_94 N_VDD_c_119_p N_C_c_196_n 6.92542e-19
cc_95 N_VDD_c_75_n N_C_c_197_n 4.58746e-19
cc_96 N_VDD_c_83_n N_C_c_197_n 8.66889e-19
cc_97 N_VDD_c_83_n N_C_c_198_n 2.22969e-19
cc_98 N_VDD_c_85_n N_C_c_198_n 2.64043e-19
cc_99 N_VDD_c_119_p N_C_c_198_n 4.74797e-19
cc_100 N_VDD_XI20.X0_PGD N_B_XI24.X0_PGS 0.00135245f
cc_101 N_VDD_XI22.X0_PGD N_B_XI24.X0_PGS 4.12959e-19
cc_102 N_VDD_c_68_n N_B_XI23.X0_PGS 0.00108553f
cc_103 N_VDD_c_68_n N_B_c_240_n 0.00256877f
cc_104 N_VDD_c_129_p N_B_c_240_n 4.12959e-19
cc_105 N_VDD_c_130_p N_B_c_242_n 0.00495207f
cc_106 N_VDD_c_89_n N_B_c_242_n 4.60491e-19
cc_107 N_VDD_XI22.X0_PGD N_A_XI23.X0_CG 4.83278e-19
cc_108 N_VDD_XI21.X0_PGD N_A_XI25.X0_PGS 0.00150004f
cc_109 N_VDD_c_85_n N_A_XI25.X0_PGS 2.05774e-19
cc_110 N_VDD_XI22.X0_PGD N_A_c_269_n 5.50272e-19
cc_111 N_VDD_XI21.X0_PGD N_A_c_270_n 3.23173e-19
cc_112 N_VDD_c_137_p N_A_c_270_n 0.00145458f
cc_113 N_VDD_c_129_p N_A_c_270_n 2.17009e-19
cc_114 N_Z_c_145_n N_C_c_194_n 2.87038e-19
cc_115 N_Z_c_146_n N_C_c_194_n 2.87038e-19
cc_116 N_Z_c_149_n N_C_c_194_n 7.3418e-19
cc_117 N_Z_c_172_n N_C_c_195_n 0.00103972f
cc_118 N_Z_c_149_n C 2.05514e-19
cc_119 N_Z_c_149_n N_C_c_196_n 0.00135375f
cc_120 N_Z_c_172_n N_C_c_196_n 2.38669e-19
cc_121 N_Z_c_149_n N_C_c_197_n 2.28309e-19
cc_122 N_Z_c_149_n N_B_XI24.X0_PGS 7.69255e-19
cc_123 N_Z_c_149_n N_B_XI23.X0_PGS 8.11898e-19
cc_124 N_Z_c_149_n N_B_c_234_n 2.98201e-19
cc_125 N_Z_c_149_n N_B_c_242_n 2.18216e-19
cc_126 N_Z_c_149_n N_A_XI23.X0_CG 7.49661e-19
cc_127 N_Z_c_149_n N_A_c_274_n 2.18216e-19
cc_128 N_Z_c_149_n N_A_c_259_n 2.14102e-19
cc_129 N_Z_c_149_n N_A_c_261_n 2.49841e-19
cc_130 N_Z_c_151_n N_A_c_261_n 4.09814e-19
cc_131 N_C_c_194_n N_B_XI24.X0_PGS 0.00849032f
cc_132 N_C_c_197_n N_B_XI24.X0_PGS 3.76133e-19
cc_133 N_C_c_194_n N_B_XI23.X0_PGS 6.67601e-19
cc_134 N_C_c_195_n N_B_XI23.X0_PGS 4.29907e-19
cc_135 N_C_c_195_n N_A_XI23.X0_CG 0.00200107f
cc_136 N_C_c_195_n N_A_XI25.X0_PGS 0.00801113f
cc_137 N_C_c_196_n N_A_c_261_n 0.00114292f
cc_138 N_B_XI24.X0_PGS N_A_XI23.X0_CG 8.40291e-19
cc_139 N_B_XI23.X0_PGS N_A_XI23.X0_CG 0.00774979f
cc_140 N_B_c_234_n N_A_c_259_n 3.39698e-19
cc_141 N_B_c_242_n N_A_c_259_n 3.48267e-19
cc_142 N_B_c_234_n N_A_c_269_n 3.48267e-19
cc_143 N_B_c_242_n N_A_c_269_n 5.15124e-19
*
.ends
*
*
.subckt MIN3_HPNW12 A B C Y VDD VSS
xgate (VSS VDD Y C B A) G3_MIN3_T6_N3
.ends
*
* File: G4_MUX2_N3.pex.netlist
* Created: Tue Mar 15 11:34:09 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_MUX2_N3_VDD 2 4 6 8 10 12 14 16 18 20 38 49 51 58 64 72 77 81 84
+ 85 89 93 95 96 99 101 105 107 111 113 115 120 122 124 125 126 127 128 134 139
+ 148 Vss
c131 148 Vss 0.00702165f
c132 139 Vss 0.00462928f
c133 134 Vss 0.00483792f
c134 128 Vss 4.52364e-19
c135 127 Vss 2.39889e-19
c136 126 Vss 4.24532e-19
c137 125 Vss 2.39889e-19
c138 122 Vss 0.00282332f
c139 120 Vss 0.0106931f
c140 115 Vss 0.00186946f
c141 113 Vss 0.006422f
c142 111 Vss 8.80889e-19
c143 107 Vss 0.00804399f
c144 105 Vss 0.00134677f
c145 101 Vss 0.00193004f
c146 99 Vss 3.98903e-19
c147 96 Vss 6.1175e-19
c148 95 Vss 0.00358057f
c149 93 Vss 0.00108621f
c150 89 Vss 0.00158874f
c151 86 Vss 0.00176185f
c152 85 Vss 0.0067647f
c153 84 Vss 0.00573691f
c154 81 Vss 0.00850511f
c155 77 Vss 0.00688835f
c156 72 Vss 0.00820121f
c157 64 Vss 8.40042e-20
c158 59 Vss 0.0806024f
c159 58 Vss 0.103898f
c160 49 Vss 0.0356247f
c161 48 Vss 0.101315f
c162 39 Vss 0.0367394f
c163 38 Vss 0.101469f
c164 18 Vss 0.188795f
c165 16 Vss 0.00143493f
c166 14 Vss 0.191141f
c167 10 Vss 0.187414f
c168 8 Vss 0.189706f
c169 6 Vss 0.190935f
c170 4 Vss 0.189249f
r171 121 128 0.551426
r172 121 122 5.50157
r173 120 128 0.551426
r174 119 120 18.3386
r175 115 128 0.0828784
r176 115 117 1.82344
r177 114 127 0.494161
r178 113 119 0.652036
r179 113 114 10.1279
r180 111 148 1.16709
r181 109 127 0.128424
r182 109 111 2.16729
r183 108 126 0.494161
r184 107 122 0.652036
r185 107 108 13.0037
r186 103 126 0.128424
r187 103 105 6.16843
r188 102 125 0.494161
r189 101 127 0.494161
r190 101 102 4.58464
r191 99 139 1.16709
r192 97 125 0.128424
r193 97 99 2.16729
r194 95 126 0.494161
r195 95 96 7.46046
r196 93 134 1.16709
r197 91 96 0.652036
r198 91 93 2.16729
r199 87 124 0.306046
r200 87 89 1.82344
r201 85 125 0.494161
r202 85 86 10.1279
r203 84 124 0.349767
r204 83 86 0.652036
r205 83 84 5.50157
r206 81 117 1.16709
r207 77 105 1.16709
r208 72 89 1.16709
r209 64 148 0.0476429
r210 64 66 1.92555
r211 59 66 0.5835
r212 58 60 0.652036
r213 58 59 2.8008
r214 55 66 0.0685365
r215 51 139 0.0476429
r216 49 51 1.45875
r217 48 52 0.652036
r218 48 51 1.45875
r219 45 49 0.652036
r220 41 134 0.0476429
r221 39 41 1.45875
r222 38 42 0.652036
r223 38 41 1.45875
r224 35 39 0.652036
r225 20 81 0.123773
r226 18 60 5.1348
r227 16 77 0.123773
r228 14 55 5.1348
r229 12 77 0.123773
r230 10 52 5.1348
r231 8 45 5.1348
r232 6 35 5.1348
r233 4 42 5.1348
r234 2 72 0.123773
.ends

.subckt PM_G4_MUX2_N3_VSS 2 4 6 8 10 12 14 16 18 20 38 39 41 48 49 59 72 77 81
+ 84 89 94 99 104 109 118 123 132 140 141 146 152 153 158 164 170 172 177 179
+ 181 182 183 184 185 Vss
c124 185 Vss 4.28045e-19
c125 184 Vss 3.62111e-19
c126 183 Vss 3.91906e-19
c127 182 Vss 3.21876e-19
c128 179 Vss 0.00582395f
c129 177 Vss 0.00193102f
c130 172 Vss 0.00135159f
c131 170 Vss 0.00259462f
c132 164 Vss 0.00592925f
c133 158 Vss 0.00385718f
c134 153 Vss 5.94991e-19
c135 152 Vss 0.00258264f
c136 147 Vss 0.00135554f
c137 146 Vss 0.00523922f
c138 141 Vss 0.00344346f
c139 140 Vss 0.00104615f
c140 132 Vss 0.00918942f
c141 123 Vss 0.00383026f
c142 118 Vss 0.00413434f
c143 109 Vss 3.63432e-19
c144 104 Vss 0.0017597f
c145 99 Vss 0.00131312f
c146 94 Vss 6.11605e-19
c147 89 Vss 0.00100326f
c148 84 Vss 0.00146588f
c149 81 Vss 0.00807726f
c150 77 Vss 0.00622224f
c151 72 Vss 0.0101685f
c152 65 Vss 0.0783825f
c153 59 Vss 0.0350566f
c154 58 Vss 0.0688416f
c155 49 Vss 0.0347733f
c156 48 Vss 0.100364f
c157 41 Vss 8.95828e-20
c158 39 Vss 0.0350852f
c159 38 Vss 0.0994129f
c160 20 Vss 0.190105f
c161 16 Vss 0.189529f
c162 14 Vss 0.00143493f
c163 12 Vss 0.189243f
c164 10 Vss 0.189689f
c165 4 Vss 0.190073f
c166 2 Vss 0.189016f
r167 178 185 0.551426
r168 178 179 18.3386
r169 177 185 0.551426
r170 176 177 5.50157
r171 172 185 0.0828784
r172 171 184 0.494161
r173 170 179 0.652036
r174 170 171 4.41793
r175 166 184 0.128424
r176 165 183 0.494161
r177 164 176 0.652036
r178 164 165 13.0037
r179 160 183 0.128424
r180 159 182 0.494161
r181 158 184 0.494161
r182 158 159 10.2946
r183 154 182 0.128424
r184 152 183 0.494161
r185 152 153 7.46046
r186 148 153 0.652036
r187 146 182 0.494161
r188 146 147 10.1279
r189 142 181 0.306046
r190 141 147 0.652036
r191 140 181 0.349767
r192 140 141 5.50157
r193 109 172 1.82344
r194 104 132 1.16709
r195 104 166 2.16729
r196 99 160 6.16843
r197 94 123 1.16709
r198 94 154 2.16729
r199 89 118 1.16709
r200 89 148 2.16729
r201 84 142 1.82344
r202 81 109 1.16709
r203 77 99 1.16709
r204 72 84 1.16709
r205 65 132 0.0476429
r206 63 65 1.8672
r207 60 63 0.0685365
r208 58 63 0.5835
r209 58 59 2.8008
r210 55 59 0.652036
r211 51 123 0.0476429
r212 49 51 1.45875
r213 48 52 0.652036
r214 48 51 1.45875
r215 45 49 0.652036
r216 41 118 0.0476429
r217 39 41 1.45875
r218 38 42 0.652036
r219 38 41 1.45875
r220 35 39 0.652036
r221 20 60 5.1348
r222 18 81 0.123773
r223 16 55 5.1348
r224 14 77 0.123773
r225 12 52 5.1348
r226 10 45 5.1348
r227 8 77 0.123773
r228 6 72 0.123773
r229 4 35 5.1348
r230 2 42 5.1348
.ends

.subckt PM_G4_MUX2_N3_ZI 2 4 6 8 10 12 27 28 43 47 50 55 60 65 81 82 91 Vss
c65 82 Vss 9.82283e-19
c66 81 Vss 0.00344769f
c67 65 Vss 0.00531208f
c68 60 Vss 0.00107621f
c69 55 Vss 0.00120586f
c70 50 Vss 0.00184713f
c71 47 Vss 0.00665316f
c72 43 Vss 0.00665316f
c73 28 Vss 0.206957f
c74 27 Vss 8.47557e-20
c75 23 Vss 0.0247918f
c76 12 Vss 0.00143493f
c77 10 Vss 0.00143493f
c78 4 Vss 0.189507f
c79 2 Vss 0.180667f
r80 87 91 0.494161
r81 83 91 0.494161
r82 81 91 0.128424
r83 81 82 13.2121
r84 77 82 0.652036
r85 60 87 5.50157
r86 55 83 6.16843
r87 50 65 1.16709
r88 50 77 2.16729
r89 47 60 1.16709
r90 43 55 1.16709
r91 31 65 0.0476429
r92 29 31 0.326018
r93 29 31 0.1167
r94 28 32 0.652036
r95 28 31 6.7686
r96 27 65 0.357321
r97 23 31 0.326018
r98 23 27 0.40845
r99 12 47 0.123773
r100 10 43 0.123773
r101 8 47 0.123773
r102 6 43 0.123773
r103 4 32 5.1348
r104 2 27 4.72635
.ends

.subckt PM_G4_MUX2_N3_Z 2 4 13 16 Vss
c13 16 Vss 2.03714e-19
c14 13 Vss 0.00452755f
c15 4 Vss 0.00143493f
r16 16 19 0.0416786
r17 13 19 1.16709
r18 4 13 0.123773
r19 2 13 0.123773
.ends

.subckt PM_G4_MUX2_N3_SELI 2 4 6 8 18 21 29 33 36 38 43 44 52 57 71 76 77 Vss
c72 77 Vss 8.29462e-19
c73 76 Vss 1.71087e-19
c74 71 Vss 0.00163664f
c75 57 Vss 0.00292618f
c76 52 Vss 0.00318194f
c77 44 Vss 0.00264419f
c78 43 Vss 8.75265e-19
c79 38 Vss 0.00210957f
c80 36 Vss 3.78531e-19
c81 33 Vss 0.00302148f
c82 29 Vss 0.00524134f
c83 21 Vss 0.16662f
c84 18 Vss 7.81442e-20
c85 6 Vss 0.166657f
c86 4 Vss 0.00143493f
r87 76 77 0.655813
r88 75 76 3.501
r89 71 75 0.655813
r90 43 52 1.16709
r91 43 71 2.00578
r92 43 44 0.513084
r93 38 57 1.16709
r94 38 77 2.00578
r95 36 44 7.46046
r96 31 36 0.652036
r97 31 33 7.91893
r98 29 33 1.16709
r99 21 57 0.50025
r100 18 52 0.50025
r101 8 21 4.37625
r102 6 18 4.37625
r103 4 29 0.123773
r104 2 29 0.123773
.ends

.subckt PM_G4_MUX2_N3_SEL 2 4 6 8 16 17 22 26 33 36 40 41 44 45 47 49 56 57 59
+ 64 69 Vss
c65 69 Vss 0.00293892f
c66 64 Vss 0.00330355f
c67 59 Vss 0.00281287f
c68 57 Vss 3.29949e-19
c69 56 Vss 0.00195862f
c70 49 Vss 4.84367e-19
c71 47 Vss 0.00164668f
c72 45 Vss 5.48919e-19
c73 44 Vss 0.00192809f
c74 41 Vss 0.00187197f
c75 36 Vss 8.44333e-20
c76 33 Vss 9.14819e-20
c77 26 Vss 0.16662f
c78 22 Vss 0.180313f
c79 20 Vss 0.0247918f
c80 17 Vss 0.0358843f
c81 16 Vss 0.179072f
c82 8 Vss 0.16662f
c83 2 Vss 0.193774f
r84 55 64 1.16709
r85 55 57 0.4602
r86 55 56 0.52504
r87 52 59 1.16709
r88 49 52 0.5835
r89 47 69 1.16709
r90 45 47 2.00578
r91 43 45 0.655813
r92 43 44 3.501
r93 41 44 0.655813
r94 41 57 1.49522
r95 40 56 2.58407
r96 38 49 0.0685365
r97 38 40 2.00057
r98 36 59 0.0476429
r99 33 69 0.50025
r100 26 64 0.50025
r101 22 59 0.357321
r102 20 36 0.326018
r103 20 22 0.40845
r104 17 36 6.7686
r105 16 36 0.326018
r106 16 36 0.1167
r107 13 17 0.652036
r108 8 33 4.37625
r109 6 26 4.37625
r110 4 22 4.72635
r111 2 13 5.1348
.ends

.subckt PM_G4_MUX2_N3_B 2 4 14 17 20 23 Vss
c30 23 Vss 0.00439028f
c31 20 Vss 2.87096e-19
c32 14 Vss 0.0853197f
c33 2 Vss 0.656289f
r34 20 23 1.16709
r35 17 20 0.109406
r36 14 23 0.0476429
r37 11 14 1.92555
r38 7 11 0.0685365
r39 4 7 5.1348
r40 2 4 17.9718
.ends

.subckt PM_G4_MUX2_N3_A 2 4 12 14 20 23 Vss
c24 23 Vss 0.00548676f
c25 20 Vss 2.95003e-19
c26 14 Vss 0.0835366f
c27 12 Vss 8.63834e-20
c28 2 Vss 0.664171f
r29 17 23 1.16709
r30 17 20 0.0364688
r31 12 23 0.0476429
r32 12 14 1.92555
r33 7 14 0.0685365
r34 2 4 17.9718
r35 2 7 5.1348
.ends

.subckt G4_MUX2_N3  VDD VSS Z SEL B A
*
* A	A
* B	B
* SEL	SEL
* Z	Z
* VSS	VSS
* VDD	VDD
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_ZI_XI6.X0_CG N_VSS_XI6.X0_PGS
+ N_VDD_XI6.X0_S TIGFET_HPNW12
XI12.X0 N_SELI_XI12.X0_D N_VDD_XI12.X0_PGD N_SEL_XI12.X0_CG N_VDD_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW12
XI5.X0 N_Z_XI5.X0_D N_VDD_XI5.X0_PGD N_ZI_XI5.X0_CG N_VDD_XI5.X0_PGS
+ N_VSS_XI5.X0_S TIGFET_HPNW12
XI13.X0 N_SELI_XI13.X0_D N_VSS_XI13.X0_PGD N_SEL_XI13.X0_CG N_VSS_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW12
XI17.X0 N_ZI_XI17.X0_D N_VDD_XI17.X0_PGD N_SELI_XI17.X0_CG N_B_XI17.X0_PGS
+ N_VSS_XI17.X0_S TIGFET_HPNW12
XI15.X0 N_ZI_XI15.X0_D N_VSS_XI15.X0_PGD N_SEL_XI15.X0_CG N_B_XI15.X0_PGS
+ N_VDD_XI15.X0_S TIGFET_HPNW12
XI16.X0 N_ZI_XI16.X0_D N_VDD_XI16.X0_PGD N_SEL_XI16.X0_CG N_A_XI16.X0_PGS
+ N_VSS_XI16.X0_S TIGFET_HPNW12
XI14.X0 N_ZI_XI14.X0_D N_VSS_XI14.X0_PGD N_SELI_XI14.X0_CG N_A_XI14.X0_PGS
+ N_VDD_XI14.X0_S TIGFET_HPNW12
*
x_PM_G4_MUX2_N3_VDD N_VDD_XI6.X0_S N_VDD_XI12.X0_PGD N_VDD_XI12.X0_PGS
+ N_VDD_XI5.X0_PGD N_VDD_XI5.X0_PGS N_VDD_XI13.X0_S N_VDD_XI17.X0_PGD
+ N_VDD_XI15.X0_S N_VDD_XI16.X0_PGD N_VDD_XI14.X0_S N_VDD_c_12_p N_VDD_c_8_p
+ N_VDD_c_102_p N_VDD_c_127_p N_VDD_c_92_p N_VDD_c_86_p N_VDD_c_15_p
+ N_VDD_c_74_p N_VDD_c_10_p N_VDD_c_9_p N_VDD_c_17_p N_VDD_c_22_p N_VDD_c_13_p
+ N_VDD_c_49_p N_VDD_c_20_p N_VDD_c_16_p N_VDD_c_5_p N_VDD_c_14_p N_VDD_c_29_p
+ N_VDD_c_34_p N_VDD_c_61_p N_VDD_c_30_p N_VDD_c_33_p VDD N_VDD_c_52_p
+ N_VDD_c_56_p N_VDD_c_59_p N_VDD_c_66_p N_VDD_c_25_p N_VDD_c_21_p N_VDD_c_100_p
+ Vss PM_G4_MUX2_N3_VDD
x_PM_G4_MUX2_N3_VSS N_VSS_XI6.X0_PGD N_VSS_XI6.X0_PGS N_VSS_XI12.X0_S
+ N_VSS_XI5.X0_S N_VSS_XI13.X0_PGD N_VSS_XI13.X0_PGS N_VSS_XI17.X0_S
+ N_VSS_XI15.X0_PGD N_VSS_XI16.X0_S N_VSS_XI14.X0_PGD N_VSS_c_139_n
+ N_VSS_c_141_n N_VSS_c_202_p N_VSS_c_246_p N_VSS_c_143_n N_VSS_c_145_n
+ N_VSS_c_226_p N_VSS_c_146_n N_VSS_c_205_p N_VSS_c_148_n N_VSS_c_149_n
+ N_VSS_c_153_n N_VSS_c_157_n N_VSS_c_162_n N_VSS_c_165_n N_VSS_c_167_n
+ N_VSS_c_170_n N_VSS_c_174_n N_VSS_c_176_n N_VSS_c_177_n N_VSS_c_179_n
+ N_VSS_c_181_n N_VSS_c_184_n N_VSS_c_185_n N_VSS_c_188_n N_VSS_c_191_n
+ N_VSS_c_192_n N_VSS_c_193_n N_VSS_c_194_n VSS N_VSS_c_198_n N_VSS_c_199_n
+ N_VSS_c_200_n N_VSS_c_201_n Vss PM_G4_MUX2_N3_VSS
x_PM_G4_MUX2_N3_ZI N_ZI_XI6.X0_CG N_ZI_XI5.X0_CG N_ZI_XI17.X0_D N_ZI_XI15.X0_D
+ N_ZI_XI16.X0_D N_ZI_XI14.X0_D N_ZI_c_271_n N_ZI_c_256_n N_ZI_c_257_n
+ N_ZI_c_258_n N_ZI_c_276_n N_ZI_c_262_n N_ZI_c_264_n N_ZI_c_296_p N_ZI_c_270_n
+ N_ZI_c_290_n N_ZI_c_306_p Vss PM_G4_MUX2_N3_ZI
x_PM_G4_MUX2_N3_Z N_Z_XI6.X0_D N_Z_XI5.X0_D N_Z_c_321_n Z Vss PM_G4_MUX2_N3_Z
x_PM_G4_MUX2_N3_SELI N_SELI_XI12.X0_D N_SELI_XI13.X0_D N_SELI_XI17.X0_CG
+ N_SELI_XI14.X0_CG N_SELI_c_334_n N_SELI_c_404_p N_SELI_c_335_n N_SELI_c_338_n
+ N_SELI_c_361_n N_SELI_c_341_n N_SELI_c_342_n N_SELI_c_343_n N_SELI_c_346_n
+ N_SELI_c_347_n N_SELI_c_357_n N_SELI_c_371_n N_SELI_c_374_n Vss
+ PM_G4_MUX2_N3_SELI
x_PM_G4_MUX2_N3_SEL N_SEL_XI12.X0_CG N_SEL_XI13.X0_CG N_SEL_XI15.X0_CG
+ N_SEL_XI16.X0_CG N_SEL_c_406_n N_SEL_c_422_n N_SEL_c_456_p N_SEL_c_457_p
+ N_SEL_c_467_p N_SEL_c_415_n SEL N_SEL_c_407_n N_SEL_c_408_n N_SEL_c_429_n
+ N_SEL_c_409_n N_SEL_c_418_n N_SEL_c_411_n N_SEL_c_445_n N_SEL_c_420_n
+ N_SEL_c_448_n N_SEL_c_413_n Vss PM_G4_MUX2_N3_SEL
x_PM_G4_MUX2_N3_B N_B_XI17.X0_PGS N_B_XI15.X0_PGS N_B_c_477_n B N_B_c_471_n
+ N_B_c_473_n Vss PM_G4_MUX2_N3_B
x_PM_G4_MUX2_N3_A N_A_XI16.X0_PGS N_A_XI14.X0_PGS N_A_c_520_n N_A_c_503_n A
+ N_A_c_509_n Vss PM_G4_MUX2_N3_A
cc_1 N_VDD_XI5.X0_PGD N_VSS_XI6.X0_PGD 0.00200866f
cc_2 N_VDD_XI12.X0_PGS N_VSS_XI6.X0_PGS 2.44446e-19
cc_3 N_VDD_XI12.X0_PGD N_VSS_XI13.X0_PGD 0.00195824f
cc_4 N_VDD_XI5.X0_PGS N_VSS_XI13.X0_PGS 2.27381e-19
cc_5 N_VDD_c_5_p N_VSS_XI13.X0_PGS 2.10824e-19
cc_6 N_VDD_XI17.X0_PGD N_VSS_XI15.X0_PGD 2.31533e-19
cc_7 N_VDD_XI16.X0_PGD N_VSS_XI14.X0_PGD 2.31533e-19
cc_8 N_VDD_c_8_p N_VSS_c_139_n 0.00200866f
cc_9 N_VDD_c_9_p N_VSS_c_139_n 3.89167e-19
cc_10 N_VDD_c_10_p N_VSS_c_141_n 4.28478e-19
cc_11 N_VDD_c_9_p N_VSS_c_141_n 4.0633e-19
cc_12 N_VDD_c_12_p N_VSS_c_143_n 0.00195824f
cc_13 N_VDD_c_13_p N_VSS_c_143_n 3.10186e-19
cc_14 N_VDD_c_14_p N_VSS_c_145_n 9.06483e-19
cc_15 N_VDD_c_15_p N_VSS_c_146_n 3.23931e-19
cc_16 N_VDD_c_16_p N_VSS_c_146_n 2.74986e-19
cc_17 N_VDD_c_17_p N_VSS_c_148_n 4.89302e-19
cc_18 N_VDD_c_10_p N_VSS_c_149_n 8.67538e-19
cc_19 N_VDD_c_9_p N_VSS_c_149_n 0.00141228f
cc_20 N_VDD_c_20_p N_VSS_c_149_n 8.83788e-19
cc_21 N_VDD_c_21_p N_VSS_c_149_n 3.48267e-19
cc_22 N_VDD_c_22_p N_VSS_c_153_n 8.50587e-19
cc_23 N_VDD_c_13_p N_VSS_c_153_n 0.00141228f
cc_24 N_VDD_c_5_p N_VSS_c_153_n 0.00180638f
cc_25 N_VDD_c_25_p N_VSS_c_153_n 3.48267e-19
cc_26 N_VDD_c_10_p N_VSS_c_157_n 2.85826e-19
cc_27 N_VDD_c_20_p N_VSS_c_157_n 3.92901e-19
cc_28 N_VDD_c_16_p N_VSS_c_157_n 2.9533e-19
cc_29 N_VDD_c_29_p N_VSS_c_157_n 7.06793e-19
cc_30 N_VDD_c_30_p N_VSS_c_157_n 4.71075e-19
cc_31 N_VDD_c_5_p N_VSS_c_162_n 2.93442e-19
cc_32 N_VDD_c_14_p N_VSS_c_162_n 0.00161703f
cc_33 N_VDD_c_33_p N_VSS_c_162_n 4.28751e-19
cc_34 N_VDD_c_34_p N_VSS_c_165_n 3.5277e-19
cc_35 N_VDD_c_30_p N_VSS_c_165_n 0.00187494f
cc_36 N_VDD_c_10_p N_VSS_c_167_n 3.66936e-19
cc_37 N_VDD_c_9_p N_VSS_c_167_n 0.00114511f
cc_38 N_VDD_c_21_p N_VSS_c_167_n 6.489e-19
cc_39 N_VDD_c_22_p N_VSS_c_170_n 3.82294e-19
cc_40 N_VDD_c_13_p N_VSS_c_170_n 0.00114511f
cc_41 N_VDD_c_5_p N_VSS_c_170_n 9.55349e-19
cc_42 N_VDD_c_25_p N_VSS_c_170_n 6.46219e-19
cc_43 N_VDD_c_14_p N_VSS_c_174_n 2.26455e-19
cc_44 N_VDD_c_33_p N_VSS_c_174_n 5.86293e-19
cc_45 N_VDD_c_10_p N_VSS_c_176_n 3.30364e-19
cc_46 N_VDD_c_22_p N_VSS_c_177_n 3.85245e-19
cc_47 N_VDD_c_5_p N_VSS_c_177_n 2.91233e-19
cc_48 N_VDD_c_13_p N_VSS_c_179_n 0.00427835f
cc_49 N_VDD_c_49_p N_VSS_c_179_n 0.00166784f
cc_50 N_VDD_c_9_p N_VSS_c_181_n 0.00425881f
cc_51 N_VDD_c_16_p N_VSS_c_181_n 0.00135965f
cc_52 N_VDD_c_52_p N_VSS_c_181_n 0.0010575f
cc_53 N_VDD_c_9_p N_VSS_c_184_n 0.00176255f
cc_54 N_VDD_c_13_p N_VSS_c_185_n 0.00138037f
cc_55 N_VDD_c_14_p N_VSS_c_185_n 0.00614137f
cc_56 N_VDD_c_56_p N_VSS_c_185_n 0.00120833f
cc_57 N_VDD_c_16_p N_VSS_c_188_n 0.00135965f
cc_58 N_VDD_c_34_p N_VSS_c_188_n 0.00823017f
cc_59 N_VDD_c_59_p N_VSS_c_188_n 0.00103007f
cc_60 N_VDD_c_14_p N_VSS_c_191_n 0.00457914f
cc_61 N_VDD_c_61_p N_VSS_c_192_n 4.01154e-19
cc_62 N_VDD_c_30_p N_VSS_c_193_n 0.0041789f
cc_63 N_VDD_c_5_p N_VSS_c_194_n 4.46614e-19
cc_64 N_VDD_c_30_p N_VSS_c_194_n 0.00867926f
cc_65 N_VDD_c_33_p N_VSS_c_194_n 0.00355235f
cc_66 N_VDD_c_66_p N_VSS_c_194_n 0.0010706f
cc_67 N_VDD_c_13_p N_VSS_c_198_n 7.23159e-19
cc_68 N_VDD_c_16_p N_VSS_c_199_n 0.00111918f
cc_69 N_VDD_c_14_p N_VSS_c_200_n 7.61747e-19
cc_70 N_VDD_c_30_p N_VSS_c_201_n 9.16632e-19
cc_71 N_VDD_XI5.X0_PGD N_ZI_c_256_n 3.96029e-19
cc_72 N_VDD_c_34_p N_ZI_c_257_n 2.74986e-19
cc_73 N_VDD_c_15_p N_ZI_c_258_n 3.43419e-19
cc_74 N_VDD_c_74_p N_ZI_c_258_n 3.43419e-19
cc_75 N_VDD_c_5_p N_ZI_c_258_n 3.48267e-19
cc_76 N_VDD_c_61_p N_ZI_c_258_n 3.72199e-19
cc_77 N_VDD_c_34_p N_ZI_c_262_n 2.9533e-19
cc_78 N_VDD_c_30_p N_ZI_c_262_n 9.20678e-19
cc_79 N_VDD_c_15_p N_ZI_c_264_n 3.48267e-19
cc_80 N_VDD_c_74_p N_ZI_c_264_n 3.48267e-19
cc_81 N_VDD_c_5_p N_ZI_c_264_n 4.99861e-19
cc_82 N_VDD_c_14_p N_ZI_c_264_n 3.21336e-19
cc_83 N_VDD_c_61_p N_ZI_c_264_n 5.226e-19
cc_84 N_VDD_c_30_p N_ZI_c_264_n 2.34601e-19
cc_85 N_VDD_c_13_p N_ZI_c_270_n 2.91231e-19
cc_86 N_VDD_c_86_p N_Z_c_321_n 3.43419e-19
cc_87 N_VDD_c_9_p N_Z_c_321_n 2.74986e-19
cc_88 N_VDD_c_17_p N_Z_c_321_n 3.72199e-19
cc_89 N_VDD_c_86_p Z 3.48267e-19
cc_90 N_VDD_c_9_p Z 3.66281e-19
cc_91 N_VDD_c_17_p Z 7.4527e-19
cc_92 N_VDD_c_92_p N_SELI_c_334_n 4.99294e-19
cc_93 N_VDD_c_15_p N_SELI_c_335_n 3.43419e-19
cc_94 N_VDD_c_13_p N_SELI_c_335_n 2.74986e-19
cc_95 N_VDD_c_5_p N_SELI_c_335_n 3.48267e-19
cc_96 N_VDD_c_15_p N_SELI_c_338_n 3.48267e-19
cc_97 N_VDD_c_13_p N_SELI_c_338_n 3.8357e-19
cc_98 N_VDD_c_5_p N_SELI_c_338_n 6.94315e-19
cc_99 N_VDD_c_30_p N_SELI_c_341_n 4.32468e-19
cc_100 N_VDD_c_100_p N_SELI_c_342_n 2.17157e-19
cc_101 N_VDD_XI5.X0_PGD N_SELI_c_343_n 2.35597e-19
cc_102 N_VDD_c_102_p N_SELI_c_343_n 2.28823e-19
cc_103 N_VDD_c_20_p N_SELI_c_343_n 2.91405e-19
cc_104 N_VDD_c_29_p N_SELI_c_346_n 2.28697e-19
cc_105 N_VDD_c_30_p N_SELI_c_347_n 3.66936e-19
cc_106 N_VDD_XI12.X0_PGD N_SEL_c_406_n 4.09718e-19
cc_107 N_VDD_c_14_p N_SEL_c_407_n 3.4535e-19
cc_108 N_VDD_c_30_p N_SEL_c_408_n 5.4414e-19
cc_109 N_VDD_c_34_p N_SEL_c_409_n 3.57377e-19
cc_110 N_VDD_c_30_p N_SEL_c_409_n 5.05119e-19
cc_111 N_VDD_c_15_p N_SEL_c_411_n 4.75243e-19
cc_112 N_VDD_c_5_p N_SEL_c_411_n 7.80048e-19
cc_113 N_VDD_c_30_p N_SEL_c_413_n 3.66936e-19
cc_114 N_VDD_c_5_p N_B_c_471_n 0.00142218f
cc_115 N_VDD_c_14_p N_B_c_471_n 0.00141439f
cc_116 N_VDD_c_5_p N_B_c_473_n 9.67317e-19
cc_117 N_VDD_c_14_p N_B_c_473_n 0.00120343f
cc_118 N_VDD_XI16.X0_PGD N_A_XI16.X0_PGS 0.00146246f
cc_119 N_VDD_c_30_p N_A_XI16.X0_PGS 0.00124298f
cc_120 N_VDD_c_34_p N_A_c_503_n 3.5103e-19
cc_121 N_VDD_c_30_p N_A_c_503_n 3.92527e-19
cc_122 N_VDD_c_29_p A 5.27373e-19
cc_123 N_VDD_c_34_p A 0.00141439f
cc_124 N_VDD_c_30_p A 5.12828e-19
cc_125 N_VDD_c_100_p A 3.44698e-19
cc_126 N_VDD_XI16.X0_PGD N_A_c_509_n 3.32271e-19
cc_127 N_VDD_c_127_p N_A_c_509_n 0.00480616f
cc_128 N_VDD_c_29_p N_A_c_509_n 3.95721e-19
cc_129 N_VDD_c_34_p N_A_c_509_n 0.00120343f
cc_130 N_VDD_c_30_p N_A_c_509_n 3.70842e-19
cc_131 N_VDD_c_100_p N_A_c_509_n 6.02643e-19
cc_132 N_VSS_c_202_p N_ZI_c_271_n 5.35095e-19
cc_133 N_VSS_XI6.X0_PGD N_ZI_c_256_n 4.09718e-19
cc_134 N_VSS_c_146_n N_ZI_c_257_n 3.43419e-19
cc_135 N_VSS_c_205_p N_ZI_c_257_n 3.43419e-19
cc_136 N_VSS_c_165_n N_ZI_c_257_n 3.48267e-19
cc_137 N_VSS_c_149_n N_ZI_c_276_n 3.27284e-19
cc_138 N_VSS_c_167_n N_ZI_c_276_n 2.15082e-19
cc_139 N_VSS_c_146_n N_ZI_c_262_n 3.48267e-19
cc_140 N_VSS_c_205_p N_ZI_c_262_n 3.48267e-19
cc_141 N_VSS_c_157_n N_ZI_c_262_n 0.00100597f
cc_142 N_VSS_c_165_n N_ZI_c_262_n 4.40384e-19
cc_143 N_VSS_c_188_n N_ZI_c_262_n 3.80707e-19
cc_144 N_VSS_c_192_n N_ZI_c_262_n 6.1924e-19
cc_145 N_VSS_c_194_n N_ZI_c_262_n 0.00228731f
cc_146 N_VSS_c_185_n N_ZI_c_264_n 3.80707e-19
cc_147 N_VSS_c_153_n N_ZI_c_270_n 2.70732e-19
cc_148 N_VSS_c_157_n N_ZI_c_270_n 4.41808e-19
cc_149 N_VSS_c_181_n N_ZI_c_270_n 7.14893e-19
cc_150 N_VSS_c_185_n N_ZI_c_270_n 0.00105381f
cc_151 N_VSS_c_179_n N_ZI_c_290_n 7.92312e-19
cc_152 N_VSS_c_146_n N_Z_c_321_n 3.43419e-19
cc_153 N_VSS_c_157_n N_Z_c_321_n 3.48267e-19
cc_154 N_VSS_c_146_n Z 3.48267e-19
cc_155 N_VSS_c_157_n Z 7.85754e-19
cc_156 N_VSS_c_226_p N_SELI_c_335_n 3.43419e-19
cc_157 N_VSS_c_148_n N_SELI_c_335_n 3.48267e-19
cc_158 N_VSS_c_226_p N_SELI_c_338_n 3.48267e-19
cc_159 N_VSS_c_148_n N_SELI_c_338_n 5.71987e-19
cc_160 N_VSS_c_194_n N_SELI_c_341_n 6.69121e-19
cc_161 N_VSS_c_146_n N_SELI_c_343_n 5.11666e-19
cc_162 N_VSS_c_157_n N_SELI_c_343_n 6.75781e-19
cc_163 N_VSS_c_181_n N_SELI_c_343_n 3.61249e-19
cc_164 N_VSS_c_174_n N_SELI_c_347_n 5.05931e-19
cc_165 N_VSS_c_188_n N_SELI_c_357_n 6.42552e-19
cc_166 N_VSS_c_194_n N_SELI_c_357_n 6.85767e-19
cc_167 N_VSS_XI13.X0_PGD N_SEL_c_406_n 4.03539e-19
cc_168 N_VSS_c_170_n N_SEL_c_415_n 5.28949e-19
cc_169 N_VSS_c_194_n N_SEL_c_408_n 2.60801e-19
cc_170 N_VSS_c_188_n N_SEL_c_409_n 2.29905e-19
cc_171 N_VSS_c_170_n N_SEL_c_418_n 2.18943e-19
cc_172 N_VSS_c_185_n N_SEL_c_411_n 3.31177e-19
cc_173 N_VSS_c_153_n N_SEL_c_420_n 2.15082e-19
cc_174 N_VSS_XI13.X0_PGS N_B_XI17.X0_PGS 0.00187616f
cc_175 N_VSS_XI15.X0_PGD N_B_XI17.X0_PGS 0.00145666f
cc_176 N_VSS_c_246_p N_B_c_477_n 0.00187616f
cc_177 N_VSS_c_162_n N_B_c_471_n 3.92469e-19
cc_178 N_VSS_c_174_n N_B_c_471_n 3.5189e-19
cc_179 N_VSS_c_185_n N_B_c_471_n 2.15119e-19
cc_180 N_VSS_XI15.X0_PGD N_B_c_473_n 3.23173e-19
cc_181 N_VSS_c_145_n N_B_c_473_n 0.00295829f
cc_182 N_VSS_c_162_n N_B_c_473_n 3.5189e-19
cc_183 N_VSS_c_170_n N_B_c_473_n 6.40394e-19
cc_184 N_VSS_c_174_n N_B_c_473_n 6.81736e-19
cc_185 N_VSS_c_188_n A 2.41977e-19
cc_186 N_ZI_c_256_n N_Z_c_321_n 6.90199e-19
cc_187 N_ZI_c_264_n N_SELI_c_338_n 9.22717e-19
cc_188 N_ZI_c_270_n N_SELI_c_338_n 0.00230161f
cc_189 N_ZI_c_256_n N_SELI_c_361_n 3.69647e-19
cc_190 N_ZI_c_276_n N_SELI_c_361_n 0.00194838f
cc_191 N_ZI_c_296_p N_SELI_c_361_n 9.76295e-19
cc_192 N_ZI_c_264_n N_SELI_c_341_n 0.00164769f
cc_193 N_ZI_c_262_n N_SELI_c_342_n 0.00166362f
cc_194 N_ZI_c_270_n N_SELI_c_342_n 0.00145462f
cc_195 N_ZI_c_256_n N_SELI_c_343_n 8.08917e-19
cc_196 N_ZI_c_270_n N_SELI_c_343_n 0.0018158f
cc_197 N_ZI_c_262_n N_SELI_c_357_n 7.72596e-19
cc_198 N_ZI_c_270_n N_SELI_c_357_n 7.93892e-19
cc_199 N_ZI_c_262_n N_SELI_c_371_n 6.01706e-19
cc_200 N_ZI_c_264_n N_SELI_c_371_n 3.05282e-19
cc_201 N_ZI_c_306_p N_SELI_c_371_n 6.45182e-19
cc_202 N_ZI_c_264_n N_SELI_c_374_n 8.28497e-19
cc_203 N_ZI_c_256_n N_SEL_c_406_n 0.0037589f
cc_204 N_ZI_c_296_p N_SEL_c_422_n 5.93636e-19
cc_205 N_ZI_c_258_n N_SEL_c_407_n 6.40197e-19
cc_206 N_ZI_c_264_n N_SEL_c_407_n 0.00209308f
cc_207 N_ZI_c_270_n N_SEL_c_407_n 8.88094e-19
cc_208 N_ZI_c_262_n N_SEL_c_408_n 9.51454e-19
cc_209 N_ZI_c_264_n N_SEL_c_408_n 4.59089e-19
cc_210 N_ZI_c_306_p N_SEL_c_408_n 0.00107464f
cc_211 N_ZI_c_257_n N_SEL_c_429_n 6.40197e-19
cc_212 N_ZI_c_262_n N_SEL_c_429_n 0.00193202f
cc_213 N_ZI_c_270_n N_SEL_c_418_n 0.0016105f
cc_214 N_ZI_c_256_n N_SEL_c_420_n 0.00117386f
cc_215 N_ZI_XI5.X0_CG N_B_XI17.X0_PGS 0.0018458f
cc_216 N_Z_c_321_n N_SELI_c_361_n 5.76103e-19
cc_217 Z N_SELI_c_361_n 8.85628e-19
cc_218 N_SELI_c_335_n N_SEL_c_406_n 6.90199e-19
cc_219 N_SELI_c_338_n N_SEL_c_406_n 8.57466e-19
cc_220 N_SELI_c_343_n N_SEL_c_406_n 2.79929e-19
cc_221 N_SELI_c_341_n N_SEL_c_407_n 0.00141479f
cc_222 N_SELI_c_347_n N_SEL_c_407_n 9.76295e-19
cc_223 N_SELI_c_338_n N_SEL_c_408_n 3.66824e-19
cc_224 N_SELI_c_342_n N_SEL_c_429_n 0.00170409f
cc_225 N_SELI_c_346_n N_SEL_c_429_n 9.29204e-19
cc_226 N_SELI_c_341_n N_SEL_c_409_n 9.15421e-19
cc_227 N_SELI_c_338_n N_SEL_c_418_n 0.00216212f
cc_228 N_SELI_c_343_n N_SEL_c_418_n 7.61998e-19
cc_229 N_SELI_c_343_n N_SEL_c_411_n 0.00193122f
cc_230 N_SELI_c_342_n N_SEL_c_445_n 0.00200661f
cc_231 N_SELI_c_338_n N_SEL_c_420_n 0.00109331f
cc_232 N_SELI_c_343_n N_SEL_c_420_n 4.73568e-19
cc_233 N_SELI_c_341_n N_SEL_c_448_n 3.48267e-19
cc_234 N_SELI_c_342_n N_SEL_c_448_n 4.95293e-19
cc_235 N_SELI_c_346_n N_SEL_c_448_n 0.00480115f
cc_236 N_SELI_c_347_n N_SEL_c_448_n 9.11855e-19
cc_237 N_SELI_c_341_n N_SEL_c_413_n 4.56568e-19
cc_238 N_SELI_c_342_n N_SEL_c_413_n 3.48267e-19
cc_239 N_SELI_c_346_n N_SEL_c_413_n 9.03632e-19
cc_240 N_SELI_c_347_n N_SEL_c_413_n 0.00245376f
cc_241 N_SELI_XI17.X0_CG N_B_XI17.X0_PGS 4.83278e-19
cc_242 N_SELI_c_338_n N_B_XI17.X0_PGS 2.54355e-19
cc_243 N_SELI_c_343_n N_B_XI17.X0_PGS 8.44835e-19
cc_244 N_SELI_c_346_n N_B_XI17.X0_PGS 0.00126314f
cc_245 N_SELI_c_404_p N_A_XI16.X0_PGS 4.99479e-19
cc_246 N_SELI_c_347_n N_A_XI16.X0_PGS 0.001089f
cc_247 N_SEL_c_456_p N_B_XI17.X0_PGS 2.07014e-19
cc_248 N_SEL_c_457_p N_B_XI17.X0_PGS 4.77845e-19
cc_249 N_SEL_c_411_n N_B_XI17.X0_PGS 7.43585e-19
cc_250 N_SEL_c_420_n N_B_XI17.X0_PGS 0.00100354f
cc_251 N_SEL_c_448_n N_B_XI17.X0_PGS 0.00142122f
cc_252 N_SEL_c_445_n N_B_c_471_n 2.97827e-19
cc_253 N_SEL_c_448_n N_B_c_471_n 2.15082e-19
cc_254 N_SEL_c_445_n N_B_c_473_n 2.18943e-19
cc_255 N_SEL_c_448_n N_B_c_473_n 5.28949e-19
cc_256 N_SEL_XI16.X0_CG N_A_XI16.X0_PGS 4.99479e-19
cc_257 N_SEL_c_413_n N_A_XI16.X0_PGS 0.001089f
cc_258 N_SEL_c_467_p N_A_c_520_n 5.05931e-19
cc_259 N_SEL_c_409_n A 2.92011e-19
cc_260 N_SEL_c_413_n A 2.15082e-19
cc_261 N_SEL_c_409_n N_A_c_509_n 2.15082e-19
cc_262 N_B_XI17.X0_PGS N_A_XI16.X0_PGS 0.00134425f
*
.ends
*
*
.subckt MUX2_HPNW12 A B S0 Y VDD VSS
xgate (VDD VSS Y S0 B A) G4_MUX2_N3
.ends
*
* File: G3_MUXI2_N3.pex.netlist
* Created: Wed Mar  9 15:24:03 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_MUXI2_N3_VSS 2 4 6 8 10 12 14 29 39 51 55 60 63 68 73 78 83 92 101
+ 110 115 121 127 133 135 140 142 144 145 146 147 Vss
c77 147 Vss 4.28045e-19
c78 146 Vss 3.62111e-19
c79 145 Vss 3.75522e-19
c80 142 Vss 0.00603414f
c81 140 Vss 0.00196409f
c82 135 Vss 0.00134915f
c83 133 Vss 0.00261859f
c84 128 Vss 0.00128551f
c85 127 Vss 0.00634725f
c86 121 Vss 0.00397667f
c87 115 Vss 0.00552282f
c88 111 Vss 0.00129855f
c89 110 Vss 0.00492065f
c90 101 Vss 0.00967583f
c91 92 Vss 0.00411469f
c92 83 Vss 2.01624e-19
c93 78 Vss 0.0013136f
c94 73 Vss 0.00223792f
c95 68 Vss 4.13309e-19
c96 63 Vss 0.00127305f
c97 60 Vss 0.00806368f
c98 55 Vss 0.00637385f
c99 51 Vss 0.0100822f
c100 45 Vss 0.0783825f
c101 39 Vss 0.0354115f
c102 38 Vss 0.0688416f
c103 29 Vss 0.0347733f
c104 28 Vss 0.101002f
c105 14 Vss 0.189925f
c106 10 Vss 0.190498f
c107 6 Vss 0.190106f
c108 4 Vss 0.189513f
r109 141 147 0.551426
r110 141 142 18.3386
r111 140 147 0.551426
r112 139 140 5.50157
r113 135 147 0.0828784
r114 134 146 0.494161
r115 133 142 0.652036
r116 133 134 4.41793
r117 129 146 0.128424
r118 127 139 0.652036
r119 127 128 13.0037
r120 123 128 0.652036
r121 122 145 0.494161
r122 121 146 0.494161
r123 121 122 10.2946
r124 117 145 0.128424
r125 116 144 0.326018
r126 115 145 0.494161
r127 115 116 10.1279
r128 110 144 0.326018
r129 109 111 0.655813
r130 109 110 5.50157
r131 83 135 1.82344
r132 78 101 1.16709
r133 78 129 2.16729
r134 73 123 6.16843
r135 68 92 1.16709
r136 68 117 2.16729
r137 63 111 1.82344
r138 60 83 1.16709
r139 55 73 1.16709
r140 51 63 1.16709
r141 45 101 0.0476429
r142 43 45 1.8672
r143 40 43 0.0685365
r144 38 43 0.5835
r145 38 39 2.8008
r146 35 39 0.652036
r147 31 92 0.0476429
r148 29 31 1.45875
r149 28 32 0.652036
r150 28 31 1.45875
r151 25 29 0.652036
r152 14 40 5.1348
r153 12 60 0.123773
r154 10 35 5.1348
r155 8 55 0.123773
r156 6 32 5.1348
r157 4 25 5.1348
r158 2 51 0.123773
.ends

.subckt PM_G3_MUXI2_N3_VDD 2 4 6 8 10 12 14 28 38 44 52 56 60 62 63 66 68 72 74
+ 75 76 81 83 84 85 87 89 98 Vss
c91 98 Vss 0.0111734f
c92 89 Vss 0.00463585f
c93 85 Vss 4.52364e-19
c94 84 Vss 4.43941e-19
c95 83 Vss 0.00378478f
c96 81 Vss 0.0102529f
c97 76 Vss 0.00177107f
c98 75 Vss 6.09322e-19
c99 74 Vss 0.0063331f
c100 72 Vss 0.00100496f
c101 68 Vss 0.00791367f
c102 66 Vss 0.00123499f
c103 63 Vss 6.1175e-19
c104 62 Vss 0.00364703f
c105 60 Vss 8.24271e-19
c106 56 Vss 0.00850511f
c107 52 Vss 0.00631561f
c108 39 Vss 0.0806024f
c109 38 Vss 0.103898f
c110 29 Vss 0.0367394f
c111 28 Vss 0.101312f
c112 12 Vss 0.189418f
c113 10 Vss 0.00143493f
c114 8 Vss 0.191033f
c115 4 Vss 0.190935f
c116 2 Vss 0.189512f
r117 83 87 0.326018
r118 82 85 0.551426
r119 82 83 5.50157
r120 81 85 0.551426
r121 80 81 18.3386
r122 76 85 0.0828784
r123 76 78 1.82344
r124 74 80 0.652036
r125 74 75 10.1279
r126 72 98 1.16709
r127 70 75 0.652036
r128 70 72 2.16729
r129 69 84 0.494161
r130 68 87 0.326018
r131 68 69 13.0037
r132 64 84 0.128424
r133 64 66 6.16843
r134 62 84 0.494161
r135 62 63 7.46046
r136 60 89 1.16709
r137 58 63 0.652036
r138 58 60 2.16729
r139 56 78 1.16709
r140 52 66 1.16709
r141 44 98 0.0476429
r142 44 46 1.92555
r143 39 46 0.5835
r144 38 40 0.652036
r145 38 39 2.8008
r146 35 46 0.0685365
r147 31 89 0.0476429
r148 29 31 1.45875
r149 28 32 0.652036
r150 28 31 1.45875
r151 25 29 0.652036
r152 14 56 0.123773
r153 12 40 5.1348
r154 10 52 0.123773
r155 8 35 5.1348
r156 6 52 0.123773
r157 4 25 5.1348
r158 2 32 5.1348
.ends

.subckt PM_G3_MUXI2_N3_SELI 2 4 6 8 21 29 33 35 38 43 53 58 72 77 78 Vss
c62 78 Vss 8.12386e-19
c63 72 Vss 0.00203892f
c64 58 Vss 0.00238787f
c65 53 Vss 0.00260984f
c66 43 Vss 7.43568e-19
c67 38 Vss 0.00160083f
c68 36 Vss 0.00170119f
c69 35 Vss 0.00410624f
c70 33 Vss 0.00348196f
c71 29 Vss 0.00498872f
c72 21 Vss 0.166608f
c73 6 Vss 0.166608f
c74 4 Vss 0.00143493f
r75 77 78 0.655813
r76 76 77 3.501
r77 72 76 0.655813
r78 43 53 1.16709
r79 43 72 2.00578
r80 43 46 0.333429
r81 38 58 1.16709
r82 38 78 2.00578
r83 35 46 0.0685365
r84 35 36 7.46046
r85 31 36 0.652036
r86 31 33 7.91893
r87 29 33 1.16709
r88 21 58 0.50025
r89 18 53 0.50025
r90 8 21 4.37625
r91 6 18 4.37625
r92 4 29 0.123773
r93 2 29 0.123773
.ends

.subckt PM_G3_MUXI2_N3_SEL 2 4 6 8 16 22 26 37 40 42 46 51 58 63 68 72 77 78 Vss
c61 78 Vss 6.45399e-20
c62 77 Vss 9.69437e-20
c63 72 Vss 9.15408e-19
c64 68 Vss 0.00231917f
c65 63 Vss 0.00272254f
c66 58 Vss 0.00263414f
c67 51 Vss 5.38256e-19
c68 46 Vss 2.72603e-19
c69 42 Vss 0.00115861f
c70 37 Vss 0.00194091f
c71 26 Vss 0.166758f
c72 22 Vss 0.180313f
c73 20 Vss 0.0247918f
c74 17 Vss 0.0369697f
c75 16 Vss 0.191525f
c76 8 Vss 0.166608f
c77 2 Vss 0.193774f
r78 76 78 0.655813
r79 76 77 3.501
r80 72 77 0.655813
r81 54 63 1.16709
r82 54 72 2.00578
r83 51 54 0.5835
r84 49 58 1.16709
r85 46 49 0.5835
r86 42 68 1.16709
r87 42 78 2.00578
r88 38 46 0.0685365
r89 38 40 1.45875
r90 37 51 0.0685365
r91 37 40 3.12589
r92 36 58 0.0476429
r93 33 68 0.50025
r94 26 63 0.50025
r95 22 58 0.357321
r96 20 36 0.326018
r97 20 22 0.40845
r98 17 36 6.7686
r99 16 36 0.326018
r100 16 36 0.1167
r101 13 17 0.652036
r102 8 33 4.37625
r103 6 26 4.37625
r104 4 22 4.72635
r105 2 13 5.1348
.ends

.subckt PM_G3_MUXI2_N3_B 2 4 7 16 20 25 28 Vss
c23 28 Vss 0.00703355f
c24 25 Vss 5.28389e-19
c25 20 Vss 0.0287936f
c26 16 Vss 0.0658163f
c27 7 Vss 0.142278f
c28 4 Vss 0.40422f
c29 2 Vss 0.170892f
r30 22 28 1.16709
r31 22 25 0.0364688
r32 16 28 0.50025
r33 16 18 1.9839
r34 12 20 0.494161
r35 9 20 0.494161
r36 8 18 0.0685365
r37 7 20 0.128424
r38 7 8 4.7847
r39 4 12 12.3118
r40 2 9 4.49295
.ends

.subckt PM_G3_MUXI2_N3_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00389294f
c33 27 Vss 0.0072311f
c34 23 Vss 0.0072311f
c35 8 Vss 0.00143493f
c36 6 Vss 0.00143493f
r37 33 35 5.91836
r38 30 33 6.91864
r39 27 35 1.16709
r40 23 30 1.16709
r41 8 27 0.123773
r42 6 23 0.123773
r43 4 27 0.123773
r44 2 23 0.123773
.ends

.subckt PM_G3_MUXI2_N3_A 2 4 12 14 17 23 Vss
c24 23 Vss 0.00593108f
c25 17 Vss 2.08619e-19
c26 14 Vss 0.0835366f
c27 2 Vss 0.666088f
r28 20 23 1.16709
r29 17 20 0.0416786
r30 12 23 0.0476429
r31 12 14 1.92555
r32 7 14 0.0685365
r33 2 4 17.9718
r34 2 7 5.1348
.ends

.subckt G3_MUXI2_N3  VSS VDD SEL B Z A
*
* A	A
* Z	Z
* B	B
* SEL	SEL
* VDD	VDD
* VSS	VSS
XI12.X0 N_SELI_XI12.X0_D N_VDD_XI12.X0_PGD N_SEL_XI12.X0_CG N_VDD_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW12
XI13.X0 N_SELI_XI13.X0_D N_VSS_XI13.X0_PGD N_SEL_XI13.X0_CG N_VSS_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW12
XI17.X0 N_Z_XI17.X0_D N_VDD_XI17.X0_PGD N_SELI_XI17.X0_CG N_B_XI17.X0_PGS
+ N_VSS_XI17.X0_S TIGFET_HPNW12
XI15.X0 N_Z_XI15.X0_D N_VSS_XI15.X0_PGD N_SEL_XI15.X0_CG N_B_XI15.X0_PGS
+ N_VDD_XI15.X0_S TIGFET_HPNW12
XI16.X0 N_Z_XI16.X0_D N_VDD_XI16.X0_PGD N_SEL_XI16.X0_CG N_A_XI16.X0_PGS
+ N_VSS_XI16.X0_S TIGFET_HPNW12
XI14.X0 N_Z_XI14.X0_D N_VSS_XI14.X0_PGD N_SELI_XI14.X0_CG N_A_XI14.X0_PGS
+ N_VDD_XI14.X0_S TIGFET_HPNW12
*
x_PM_G3_MUXI2_N3_VSS N_VSS_XI12.X0_S N_VSS_XI13.X0_PGD N_VSS_XI13.X0_PGS
+ N_VSS_XI17.X0_S N_VSS_XI15.X0_PGD N_VSS_XI16.X0_S N_VSS_XI14.X0_PGD
+ N_VSS_c_4_p N_VSS_c_20_p N_VSS_c_44_p N_VSS_c_67_p N_VSS_c_69_p N_VSS_c_45_p
+ N_VSS_c_5_p N_VSS_c_26_p N_VSS_c_17_p N_VSS_c_27_p N_VSS_c_9_p N_VSS_c_19_p
+ N_VSS_c_6_p N_VSS_c_10_p N_VSS_c_11_p N_VSS_c_28_p N_VSS_c_24_p N_VSS_c_30_p
+ N_VSS_c_32_p N_VSS_c_33_p VSS N_VSS_c_12_p N_VSS_c_25_p N_VSS_c_34_p Vss
+ PM_G3_MUXI2_N3_VSS
x_PM_G3_MUXI2_N3_VDD N_VDD_XI12.X0_PGD N_VDD_XI12.X0_PGS N_VDD_XI13.X0_S
+ N_VDD_XI17.X0_PGD N_VDD_XI15.X0_S N_VDD_XI16.X0_PGD N_VDD_XI14.X0_S
+ N_VDD_c_81_n N_VDD_c_164_p N_VDD_c_128_p N_VDD_c_121_p N_VDD_c_144_p
+ N_VDD_c_82_n N_VDD_c_84_n N_VDD_c_90_n N_VDD_c_91_n N_VDD_c_97_n N_VDD_c_103_n
+ N_VDD_c_104_n N_VDD_c_106_n N_VDD_c_107_n N_VDD_c_108_n N_VDD_c_112_n
+ N_VDD_c_116_n N_VDD_c_117_n VDD N_VDD_c_118_n N_VDD_c_120_n Vss
+ PM_G3_MUXI2_N3_VDD
x_PM_G3_MUXI2_N3_SELI N_SELI_XI12.X0_D N_SELI_XI13.X0_D N_SELI_XI17.X0_CG
+ N_SELI_XI14.X0_CG N_SELI_c_229_p N_SELI_c_169_n N_SELI_c_171_n N_SELI_c_174_n
+ N_SELI_c_175_n N_SELI_c_188_n N_SELI_c_191_n N_SELI_c_178_n N_SELI_c_179_n
+ N_SELI_c_180_n N_SELI_c_211_p Vss PM_G3_MUXI2_N3_SELI
x_PM_G3_MUXI2_N3_SEL N_SEL_XI12.X0_CG N_SEL_XI13.X0_CG N_SEL_XI15.X0_CG
+ N_SEL_XI16.X0_CG N_SEL_c_231_n N_SEL_c_272_p N_SEL_c_273_p N_SEL_c_232_n SEL
+ N_SEL_c_233_n N_SEL_c_234_n N_SEL_c_257_n N_SEL_c_236_n N_SEL_c_260_n
+ N_SEL_c_246_n N_SEL_c_237_n N_SEL_c_239_n N_SEL_c_240_n Vss PM_G3_MUXI2_N3_SEL
x_PM_G3_MUXI2_N3_B N_B_XI17.X0_PGS N_B_XI15.X0_PGS N_B_c_292_n N_B_c_310_n
+ N_B_c_301_n B N_B_c_293_n Vss PM_G3_MUXI2_N3_B
x_PM_G3_MUXI2_N3_Z N_Z_XI17.X0_D N_Z_XI15.X0_D N_Z_XI16.X0_D N_Z_XI14.X0_D
+ N_Z_c_315_n N_Z_c_325_n N_Z_c_319_n Z Vss PM_G3_MUXI2_N3_Z
x_PM_G3_MUXI2_N3_A N_A_XI16.X0_PGS N_A_XI14.X0_PGS N_A_c_366_n N_A_c_350_n A
+ N_A_c_356_n Vss PM_G3_MUXI2_N3_A
cc_1 N_VSS_XI13.X0_PGD N_VDD_XI12.X0_PGD 0.00200584f
cc_2 N_VSS_XI15.X0_PGD N_VDD_XI17.X0_PGD 2.44446e-19
cc_3 N_VSS_XI14.X0_PGD N_VDD_XI16.X0_PGD 2.44446e-19
cc_4 N_VSS_c_4_p N_VDD_c_81_n 0.00200584f
cc_5 N_VSS_c_5_p N_VDD_c_82_n 9.64791e-19
cc_6 N_VSS_c_6_p N_VDD_c_82_n 4.10707e-19
cc_7 N_VSS_c_4_p N_VDD_c_84_n 3.89167e-19
cc_8 N_VSS_c_5_p N_VDD_c_84_n 0.00161703f
cc_9 N_VSS_c_9_p N_VDD_c_84_n 2.26455e-19
cc_10 N_VSS_c_10_p N_VDD_c_84_n 0.00442837f
cc_11 N_VSS_c_11_p N_VDD_c_84_n 0.00129625f
cc_12 N_VSS_c_12_p N_VDD_c_84_n 7.74609e-19
cc_13 N_VSS_c_10_p N_VDD_c_90_n 0.00157719f
cc_14 N_VSS_XI13.X0_PGS N_VDD_c_91_n 2.59535e-19
cc_15 N_VSS_XI15.X0_PGD N_VDD_c_91_n 2.19376e-19
cc_16 N_VSS_c_5_p N_VDD_c_91_n 0.00180638f
cc_17 N_VSS_c_17_p N_VDD_c_91_n 7.4365e-19
cc_18 N_VSS_c_9_p N_VDD_c_91_n 9.55109e-19
cc_19 N_VSS_c_19_p N_VDD_c_91_n 2.70301e-19
cc_20 N_VSS_c_20_p N_VDD_c_97_n 0.0011044f
cc_21 N_VSS_c_17_p N_VDD_c_97_n 0.00161703f
cc_22 N_VSS_c_19_p N_VDD_c_97_n 2.26455e-19
cc_23 N_VSS_c_11_p N_VDD_c_97_n 0.00590664f
cc_24 N_VSS_c_24_p N_VDD_c_97_n 0.0034989f
cc_25 N_VSS_c_25_p N_VDD_c_97_n 7.61747e-19
cc_26 N_VSS_c_26_p N_VDD_c_103_n 0.00121523f
cc_27 N_VSS_c_27_p N_VDD_c_104_n 3.5277e-19
cc_28 N_VSS_c_28_p N_VDD_c_104_n 0.00873112f
cc_29 N_VSS_c_28_p N_VDD_c_106_n 0.00155968f
cc_30 N_VSS_c_30_p N_VDD_c_107_n 4.01154e-19
cc_31 N_VSS_c_27_p N_VDD_c_108_n 0.00187494f
cc_32 N_VSS_c_32_p N_VDD_c_108_n 0.0041789f
cc_33 N_VSS_c_33_p N_VDD_c_108_n 0.0078367f
cc_34 N_VSS_c_34_p N_VDD_c_108_n 9.16632e-19
cc_35 N_VSS_c_17_p N_VDD_c_112_n 4.28751e-19
cc_36 N_VSS_c_19_p N_VDD_c_112_n 6.0691e-19
cc_37 N_VSS_c_24_p N_VDD_c_112_n 0.00108024f
cc_38 N_VSS_c_33_p N_VDD_c_112_n 0.00418449f
cc_39 N_VSS_c_11_p N_VDD_c_116_n 0.00121059f
cc_40 N_VSS_c_33_p N_VDD_c_117_n 0.00100712f
cc_41 N_VSS_c_5_p N_VDD_c_118_n 3.48267e-19
cc_42 N_VSS_c_9_p N_VDD_c_118_n 6.46219e-19
cc_43 N_VSS_c_26_p N_VDD_c_120_n 2.82095e-19
cc_44 N_VSS_c_44_p N_SELI_c_169_n 3.43419e-19
cc_45 N_VSS_c_45_p N_SELI_c_169_n 3.48267e-19
cc_46 N_VSS_c_44_p N_SELI_c_171_n 3.48267e-19
cc_47 N_VSS_c_45_p N_SELI_c_171_n 8.50248e-19
cc_48 N_VSS_c_10_p N_SELI_c_171_n 2.24858e-19
cc_49 N_VSS_c_26_p N_SELI_c_174_n 7.64616e-19
cc_50 N_VSS_c_17_p N_SELI_c_175_n 2.2375e-19
cc_51 N_VSS_c_19_p N_SELI_c_175_n 2.18171e-19
cc_52 N_VSS_c_33_p N_SELI_c_175_n 9.07743e-19
cc_53 N_VSS_c_17_p N_SELI_c_178_n 2.15082e-19
cc_54 N_VSS_c_28_p N_SELI_c_179_n 5.93394e-19
cc_55 N_VSS_c_33_p N_SELI_c_180_n 5.03655e-19
cc_56 N_VSS_XI13.X0_PGD N_SEL_c_231_n 4.23684e-19
cc_57 N_VSS_c_11_p N_SEL_c_232_n 4.38015e-19
cc_58 N_VSS_c_33_p N_SEL_c_233_n 7.91494e-19
cc_59 N_VSS_c_5_p N_SEL_c_234_n 2.10271e-19
cc_60 N_VSS_c_9_p N_SEL_c_234_n 2.26251e-19
cc_61 N_VSS_c_5_p N_SEL_c_236_n 2.15082e-19
cc_62 N_VSS_c_11_p N_SEL_c_237_n 7.83225e-19
cc_63 N_VSS_c_28_p N_SEL_c_237_n 2.12674e-19
cc_64 N_VSS_c_33_p N_SEL_c_239_n 4.36463e-19
cc_65 N_VSS_c_28_p N_SEL_c_240_n 7.26277e-19
cc_66 N_VSS_XI13.X0_PGS N_B_c_292_n 2.57132e-19
cc_67 N_VSS_c_67_p N_B_c_293_n 0.00132057f
cc_68 N_VSS_c_67_p N_Z_c_315_n 3.43419e-19
cc_69 N_VSS_c_69_p N_Z_c_315_n 3.43419e-19
cc_70 N_VSS_c_26_p N_Z_c_315_n 3.48267e-19
cc_71 N_VSS_c_27_p N_Z_c_315_n 3.48267e-19
cc_72 N_VSS_c_67_p N_Z_c_319_n 3.48267e-19
cc_73 N_VSS_c_69_p N_Z_c_319_n 3.48267e-19
cc_74 N_VSS_c_26_p N_Z_c_319_n 5.68482e-19
cc_75 N_VSS_c_27_p N_Z_c_319_n 5.71987e-19
cc_76 N_VSS_c_33_p N_Z_c_319_n 9.78034e-19
cc_77 N_VSS_c_28_p A 2.12185e-19
cc_78 N_VDD_c_121_p N_SELI_c_169_n 3.43419e-19
cc_79 N_VDD_c_84_n N_SELI_c_169_n 2.74986e-19
cc_80 N_VDD_c_91_n N_SELI_c_169_n 3.48267e-19
cc_81 N_VDD_c_121_p N_SELI_c_171_n 3.48267e-19
cc_82 N_VDD_c_84_n N_SELI_c_171_n 3.83029e-19
cc_83 N_VDD_c_91_n N_SELI_c_171_n 7.09569e-19
cc_84 N_VDD_c_108_n N_SELI_c_175_n 6.15494e-19
cc_85 N_VDD_c_128_p N_SELI_c_188_n 2.21762e-19
cc_86 N_VDD_c_103_n N_SELI_c_188_n 2.87975e-19
cc_87 N_VDD_c_120_n N_SELI_c_188_n 2.30774e-19
cc_88 N_VDD_c_103_n N_SELI_c_191_n 2.28697e-19
cc_89 N_VDD_c_108_n N_SELI_c_178_n 3.66936e-19
cc_90 N_VDD_XI12.X0_PGD N_SEL_c_231_n 4.31283e-19
cc_91 N_VDD_c_121_p N_SEL_c_232_n 4.75243e-19
cc_92 N_VDD_c_91_n N_SEL_c_232_n 8.22147e-19
cc_93 N_VDD_c_104_n N_SEL_c_233_n 2.47222e-19
cc_94 N_VDD_c_108_n N_SEL_c_233_n 6.15494e-19
cc_95 N_VDD_c_108_n N_SEL_c_246_n 3.66936e-19
cc_96 N_VDD_c_97_n N_SEL_c_237_n 3.65289e-19
cc_97 N_VDD_c_108_n N_SEL_c_239_n 2.2501e-19
cc_98 N_VDD_c_121_p N_B_c_292_n 2.35559e-19
cc_99 N_VDD_c_104_n N_Z_c_315_n 2.74986e-19
cc_100 N_VDD_c_121_p N_Z_c_325_n 3.43419e-19
cc_101 N_VDD_c_144_p N_Z_c_325_n 3.43419e-19
cc_102 N_VDD_c_91_n N_Z_c_325_n 3.48267e-19
cc_103 N_VDD_c_97_n N_Z_c_325_n 2.74986e-19
cc_104 N_VDD_c_107_n N_Z_c_325_n 3.72199e-19
cc_105 N_VDD_c_121_p N_Z_c_319_n 3.48267e-19
cc_106 N_VDD_c_144_p N_Z_c_319_n 3.48267e-19
cc_107 N_VDD_c_91_n N_Z_c_319_n 8.16241e-19
cc_108 N_VDD_c_97_n N_Z_c_319_n 3.83904e-19
cc_109 N_VDD_c_104_n N_Z_c_319_n 3.83904e-19
cc_110 N_VDD_c_107_n N_Z_c_319_n 8.08807e-19
cc_111 N_VDD_c_108_n N_Z_c_319_n 0.00135474f
cc_112 N_VDD_XI16.X0_PGD N_A_XI16.X0_PGS 0.00146246f
cc_113 N_VDD_c_108_n N_A_XI16.X0_PGS 0.00109285f
cc_114 N_VDD_c_104_n N_A_c_350_n 3.5103e-19
cc_115 N_VDD_c_108_n N_A_c_350_n 3.92527e-19
cc_116 N_VDD_c_103_n A 5.27373e-19
cc_117 N_VDD_c_104_n A 0.00141439f
cc_118 N_VDD_c_108_n A 5.06354e-19
cc_119 N_VDD_c_120_n A 3.44698e-19
cc_120 N_VDD_XI16.X0_PGD N_A_c_356_n 3.32271e-19
cc_121 N_VDD_c_164_p N_A_c_356_n 0.00480616f
cc_122 N_VDD_c_103_n N_A_c_356_n 3.95721e-19
cc_123 N_VDD_c_104_n N_A_c_356_n 0.00120343f
cc_124 N_VDD_c_108_n N_A_c_356_n 3.70842e-19
cc_125 N_VDD_c_120_n N_A_c_356_n 6.02643e-19
cc_126 N_SELI_c_169_n N_SEL_c_231_n 7.69306e-19
cc_127 N_SELI_c_171_n N_SEL_c_231_n 9.27181e-19
cc_128 N_SELI_c_174_n N_SEL_c_231_n 4.0622e-19
cc_129 N_SELI_c_188_n N_SEL_c_232_n 0.00290285f
cc_130 N_SELI_c_175_n N_SEL_c_233_n 0.00242961f
cc_131 N_SELI_c_178_n N_SEL_c_233_n 4.99367e-19
cc_132 N_SELI_c_171_n N_SEL_c_234_n 0.0024269f
cc_133 N_SELI_c_174_n N_SEL_c_234_n 0.00290285f
cc_134 N_SELI_c_191_n N_SEL_c_257_n 5.42085e-19
cc_135 N_SELI_c_171_n N_SEL_c_236_n 0.00100994f
cc_136 N_SELI_c_174_n N_SEL_c_236_n 5.63096e-19
cc_137 N_SELI_c_191_n N_SEL_c_260_n 0.00494389f
cc_138 N_SELI_c_178_n N_SEL_c_260_n 8.7809e-19
cc_139 N_SELI_c_191_n N_SEL_c_246_n 8.69867e-19
cc_140 N_SELI_c_178_n N_SEL_c_246_n 0.00494884f
cc_141 N_SELI_c_175_n N_SEL_c_237_n 0.00165721f
cc_142 N_SELI_c_188_n N_SEL_c_237_n 4.7869e-19
cc_143 N_SELI_c_179_n N_SEL_c_237_n 9.92651e-19
cc_144 N_SELI_c_211_p N_SEL_c_237_n 8.15293e-19
cc_145 N_SELI_c_171_n N_SEL_c_239_n 3.01017e-19
cc_146 N_SELI_c_180_n N_SEL_c_239_n 0.00144491f
cc_147 N_SELI_c_188_n N_SEL_c_240_n 0.00165436f
cc_148 N_SELI_c_179_n N_SEL_c_240_n 8.14736e-19
cc_149 N_SELI_XI17.X0_CG N_B_XI17.X0_PGS 4.31731e-19
cc_150 N_SELI_c_191_n N_B_XI17.X0_PGS 6.66106e-19
cc_151 N_SELI_c_171_n N_B_XI15.X0_PGS 2.97793e-19
cc_152 N_SELI_c_174_n N_B_XI15.X0_PGS 3.99745e-19
cc_153 N_SELI_c_191_n N_B_XI15.X0_PGS 5.45575e-19
cc_154 N_SELI_c_174_n N_B_c_292_n 4.07501e-19
cc_155 N_SELI_c_174_n N_B_c_301_n 5.40503e-19
cc_156 N_SELI_c_191_n N_B_c_301_n 0.00179467f
cc_157 N_SELI_c_174_n B 0.0012894f
cc_158 N_SELI_c_174_n N_B_c_293_n 0.00106912f
cc_159 N_SELI_c_171_n N_Z_c_319_n 0.00105053f
cc_160 N_SELI_c_175_n N_Z_c_319_n 0.00208341f
cc_161 N_SELI_c_188_n N_Z_c_319_n 0.00213869f
cc_162 N_SELI_c_229_p N_A_XI16.X0_PGS 4.87172e-19
cc_163 N_SELI_c_178_n N_A_XI16.X0_PGS 0.00276355f
cc_164 N_SEL_c_272_p N_B_XI15.X0_PGS 2.04953e-19
cc_165 N_SEL_c_273_p N_B_XI15.X0_PGS 4.65537e-19
cc_166 N_SEL_c_232_n N_B_XI15.X0_PGS 8.40923e-19
cc_167 N_SEL_c_236_n N_B_XI15.X0_PGS 0.00100354f
cc_168 N_SEL_c_260_n N_B_XI15.X0_PGS 0.00202689f
cc_169 N_SEL_c_232_n N_B_c_310_n 2.88938e-19
cc_170 N_SEL_c_236_n N_B_c_310_n 7.65159e-19
cc_171 N_SEL_c_236_n N_B_c_293_n 0.00115283f
cc_172 N_SEL_c_233_n N_Z_c_319_n 0.00189968f
cc_173 N_SEL_c_257_n N_Z_c_319_n 0.00240311f
cc_174 N_SEL_c_246_n N_Z_c_319_n 9.35582e-19
cc_175 N_SEL_c_237_n N_Z_c_319_n 9.65156e-19
cc_176 N_SEL_c_239_n N_Z_c_319_n 0.0021646f
cc_177 N_SEL_c_240_n N_Z_c_319_n 9.51045e-19
cc_178 N_SEL_XI16.X0_CG N_A_XI16.X0_PGS 4.87172e-19
cc_179 N_SEL_c_246_n N_A_XI16.X0_PGS 0.00276355f
cc_180 N_SEL_c_233_n N_A_c_366_n 2.18171e-19
cc_181 N_SEL_c_233_n A 2.78876e-19
cc_182 N_SEL_c_246_n A 2.15082e-19
cc_183 N_SEL_c_233_n N_A_c_356_n 2.30774e-19
cc_184 B N_Z_c_319_n 4.05731e-19
cc_185 N_B_XI17.X0_PGS N_A_XI16.X0_PGS 0.00134199f
*
.ends
*
*
.subckt MUXI2_HPNW12 A B S0 Y VDD VSS
xgate (VSS VDD S0 B Y A) G3_MUXI2_N3
.ends
*
* File: G2_NAND2_N3.pex.netlist
* Created: Sun Apr 10 19:03:25 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NAND2_N3_VSS 2 4 6 8 10 20 21 41 45 50 59 66 71 72 Vss
c25 72 Vss 8.04097e-19
c26 71 Vss 0.00222754f
c27 67 Vss 0.00133588f
c28 66 Vss 0.0113624f
c29 59 Vss 0.0053595f
c30 50 Vss 0.00153395f
c31 45 Vss 0.00130895f
c32 41 Vss 0.00965443f
c33 38 Vss 0.0299311f
c34 37 Vss 0.0299311f
c35 32 Vss 0.106916f
c36 27 Vss 0.0688416f
c37 21 Vss 0.0350852f
c38 20 Vss 0.0646396f
c39 10 Vss 0.190769f
c40 8 Vss 0.19123f
c41 6 Vss 0.189919f
c42 4 Vss 0.191018f
r43 71 73 0.652036
r44 71 72 4.33457
r45 64 72 0.652036
r46 64 66 12.5452
r47 63 67 0.655813
r48 63 66 6.50186
r49 50 59 1.16709
r50 50 73 2.16729
r51 45 67 1.82344
r52 41 45 1.16709
r53 33 38 0.494161
r54 32 34 0.652036
r55 32 33 2.9175
r56 29 38 0.128424
r57 28 37 0.494161
r58 27 38 0.494161
r59 27 28 2.8008
r60 24 37 0.128424
r61 23 59 0.0476429
r62 21 23 1.4004
r63 20 37 0.494161
r64 20 23 1.5171
r65 17 21 0.652036
r66 10 34 5.1348
r67 8 29 5.1348
r68 6 17 5.1348
r69 4 24 5.1348
r70 2 41 0.123773
.ends

.subckt PM_G2_NAND2_N3_VDD 2 4 6 15 17 22 27 30 31 33 35 36 37 41 46 48 51 57
+ Vss
c42 57 Vss 0.00431501f
c43 49 Vss 7.68513e-19
c44 48 Vss 0.00721617f
c45 46 Vss 0.00728738f
c46 41 Vss 0.00103469f
c47 37 Vss 0.0066476f
c48 36 Vss 8.606e-19
c49 35 Vss 0.0118736f
c50 33 Vss 0.00172072f
c51 31 Vss 7.81221e-19
c52 30 Vss 0.00275683f
c53 27 Vss 0.00946889f
c54 22 Vss 0.00810168f
c55 17 Vss 0.170588f
c56 15 Vss 0.0352333f
c57 2 Vss 0.220859f
r58 48 51 0.326018
r59 47 49 0.551426
r60 47 48 5.37654
r61 46 49 0.551426
r62 45 46 8.41907
r63 43 64 1.16709
r64 41 49 0.0828784
r65 41 43 1.53169
r66 39 57 1.16709
r67 37 45 0.655813
r68 37 39 4.0845
r69 35 51 0.326018
r70 35 36 15.3377
r71 31 33 1.82344
r72 30 36 0.652036
r73 29 31 0.655813
r74 29 30 5.50157
r75 27 64 0.15
r76 22 33 1.16709
r77 17 57 0.428786
r78 15 17 5.3682
r79 12 15 0.652036
r80 6 27 0.123773
r81 4 22 0.123773
r82 2 12 6.3018
.ends

.subckt PM_G2_NAND2_N3_A 1 2 20 23 28 33 Vss
c18 33 Vss 0.00403439f
c19 28 Vss 0.00239607f
c20 20 Vss 0.0017793f
c21 12 Vss 0.166936f
c22 1 Vss 0.171396f
r23 25 33 1.16709
r24 23 25 3.00086
r25 20 28 1.16709
r26 20 23 2.37568
r27 12 33 0.50025
r28 9 28 0.50025
r29 2 12 4.37625
r30 1 9 4.60965
.ends

.subckt PM_G2_NAND2_N3_Z 2 4 6 18 22 25 28 Vss
c26 25 Vss 0.00178689f
c27 22 Vss 0.0056591f
c28 18 Vss 0.00911019f
c29 6 Vss 0.00143493f
r30 30 39 1.16709
r31 28 30 6.54354
r32 25 28 7.12704
r33 22 39 0.15
r34 18 25 1.16709
r35 6 22 0.123773
r36 4 22 0.123773
r37 2 18 0.123773
.ends

.subckt PM_G2_NAND2_N3_B 2 3 9 10 13 19 Vss
c23 19 Vss 1.07412e-19
c24 13 Vss 0.244723f
c25 10 Vss 0.0357412f
c26 9 Vss 0.288308f
c27 2 Vss 0.328264f
r28 19 22 0.125036
r29 13 22 1.16709
r30 11 13 2.39235
r31 9 11 0.652036
r32 9 10 8.92755
r33 6 10 0.652036
r34 3 13 5.6016
r35 2 6 9.8028
.ends

.subckt G2_NAND2_N3  VSS VDD A Z B
*
* B	B
* Z	Z
* A	A
* VDD	VDD
* VSS	VSS
XI13.X0 N_Z_XI13.X0_D N_VDD_XI13.X0_PGD N_A_XI13.X0_CG N_B_XI13.X0_PGS
+ N_VSS_XI13.X0_S TIGFET_HPNW12
XI14.X0 N_Z_XI14.X0_D N_VSS_XI14.X0_PGD N_A_XI14.X0_CG N_VSS_XI14.X0_PGS
+ N_VDD_XI14.X0_S TIGFET_HPNW12
XI15.X0 N_Z_XI15.X0_D N_VSS_XI15.X0_PGD N_B_XI15.X0_CG N_VSS_XI15.X0_PGS
+ N_VDD_XI15.X0_S TIGFET_HPNW12
*
x_PM_G2_NAND2_N3_VSS N_VSS_XI13.X0_S N_VSS_XI14.X0_PGD N_VSS_XI14.X0_PGS
+ N_VSS_XI15.X0_PGD N_VSS_XI15.X0_PGS N_VSS_c_6_p N_VSS_c_7_p N_VSS_c_19_p
+ N_VSS_c_5_p N_VSS_c_2_p N_VSS_c_9_p VSS N_VSS_c_10_p N_VSS_c_11_p Vss
+ PM_G2_NAND2_N3_VSS
x_PM_G2_NAND2_N3_VDD N_VDD_XI13.X0_PGD N_VDD_XI14.X0_S N_VDD_XI15.X0_S
+ N_VDD_c_60_p N_VDD_c_50_p N_VDD_c_44_p N_VDD_c_45_p N_VDD_c_26_n N_VDD_c_29_n
+ N_VDD_c_30_n N_VDD_c_31_n N_VDD_c_36_n N_VDD_c_55_p N_VDD_c_48_p N_VDD_c_41_p
+ N_VDD_c_37_n VDD N_VDD_c_43_p Vss PM_G2_NAND2_N3_VDD
x_PM_G2_NAND2_N3_A N_A_XI13.X0_CG N_A_XI14.X0_CG N_A_c_68_n A N_A_c_74_n
+ N_A_c_70_n Vss PM_G2_NAND2_N3_A
x_PM_G2_NAND2_N3_Z N_Z_XI13.X0_D N_Z_XI14.X0_D N_Z_XI15.X0_D N_Z_c_86_n
+ N_Z_c_90_n N_Z_c_88_n Z Vss PM_G2_NAND2_N3_Z
x_PM_G2_NAND2_N3_B N_B_XI13.X0_PGS N_B_XI15.X0_CG N_B_c_112_n N_B_c_114_n
+ N_B_c_117_n B Vss PM_G2_NAND2_N3_B
cc_1 N_VSS_XI14.X0_PGS N_VDD_c_26_n 3.44373e-19
cc_2 N_VSS_c_2_p N_VDD_c_26_n 4.83895e-19
cc_3 VSS N_VDD_c_26_n 0.00361022f
cc_4 VSS N_VDD_c_29_n 0.00159527f
cc_5 N_VSS_c_5_p N_VDD_c_30_n 3.7872e-19
cc_6 N_VSS_c_6_p N_VDD_c_31_n 0.00194111f
cc_7 N_VSS_c_7_p N_VDD_c_31_n 3.76573e-19
cc_8 N_VSS_c_2_p N_VDD_c_31_n 0.00161703f
cc_9 N_VSS_c_9_p N_VDD_c_31_n 2.26455e-19
cc_10 N_VSS_c_10_p N_VDD_c_31_n 0.00519315f
cc_11 N_VSS_c_11_p N_VDD_c_36_n 0.00104854f
cc_12 N_VSS_XI15.X0_PGS N_VDD_c_37_n 4.24059e-19
cc_13 N_VSS_c_2_p N_VDD_c_37_n 5.47905e-19
cc_14 VSS N_VDD_c_37_n 2.38209e-19
cc_15 N_VSS_c_9_p N_A_c_68_n 2.354e-19
cc_16 VSS N_A_c_68_n 0.00258255f
cc_17 N_VSS_c_2_p N_A_c_70_n 2.15082e-19
cc_18 N_VSS_c_9_p N_A_c_70_n 4.9359e-19
cc_19 N_VSS_c_19_p N_Z_c_86_n 3.43419e-19
cc_20 N_VSS_c_5_p N_Z_c_86_n 3.48267e-19
cc_21 N_VSS_c_5_p N_Z_c_88_n 8.92744e-19
cc_22 VSS N_Z_c_88_n 0.0013442f
cc_23 N_VSS_XI14.X0_PGD N_B_c_112_n 7.63854e-19
cc_24 N_VSS_XI15.X0_PGD N_B_c_112_n 7.63854e-19
cc_25 N_VSS_XI14.X0_PGS N_B_c_114_n 9.45978e-19
cc_26 N_VDD_XI13.X0_PGD N_A_XI13.X0_CG 4.9269e-19
cc_27 N_VDD_c_41_p N_A_c_68_n 2.11067e-19
cc_28 N_VDD_XI13.X0_PGD N_A_c_74_n 4.86892e-19
cc_29 N_VDD_c_43_p N_A_c_74_n 5.00305e-19
cc_30 N_VDD_c_44_p N_Z_c_90_n 3.43419e-19
cc_31 N_VDD_c_45_p N_Z_c_90_n 3.43419e-19
cc_32 N_VDD_c_30_n N_Z_c_90_n 3.72199e-19
cc_33 N_VDD_c_31_n N_Z_c_90_n 2.82909e-19
cc_34 N_VDD_c_48_p N_Z_c_90_n 3.70313e-19
cc_35 N_VDD_XI13.X0_PGD N_Z_c_88_n 3.98301e-19
cc_36 N_VDD_c_50_p N_Z_c_88_n 6.23961e-19
cc_37 N_VDD_c_44_p N_Z_c_88_n 3.48267e-19
cc_38 N_VDD_c_45_p N_Z_c_88_n 3.48267e-19
cc_39 N_VDD_c_30_n N_Z_c_88_n 8.08807e-19
cc_40 N_VDD_c_31_n N_Z_c_88_n 5.69519e-19
cc_41 N_VDD_c_55_p N_Z_c_88_n 0.00170631f
cc_42 N_VDD_c_48_p N_Z_c_88_n 8.48488e-19
cc_43 N_VDD_c_41_p N_Z_c_88_n 0.00275333f
cc_44 N_VDD_c_43_p N_Z_c_88_n 9.31683e-19
cc_45 N_VDD_XI13.X0_PGD N_B_XI13.X0_PGS 0.00331576f
cc_46 N_VDD_c_60_p N_B_c_112_n 0.00812117f
cc_47 N_VDD_c_55_p N_B_c_117_n 3.69683e-19
cc_48 N_VDD_c_41_p N_B_c_117_n 6.28222e-19
cc_49 N_VDD_c_43_p N_B_c_117_n 0.00146481f
cc_50 N_VDD_c_31_n B 2.63427e-19
cc_51 N_VDD_c_55_p B 5.03854e-19
cc_52 N_VDD_c_41_p B 7.0924e-19
cc_53 N_VDD_c_43_p B 3.69683e-19
cc_54 N_A_c_68_n N_Z_c_88_n 0.00825864f
cc_55 N_A_c_74_n N_Z_c_88_n 8.85473e-19
cc_56 N_A_c_70_n N_Z_c_88_n 0.00100714f
cc_57 N_A_XI13.X0_CG N_B_XI13.X0_PGS 4.97429e-19
cc_58 N_A_c_68_n N_B_XI13.X0_PGS 5.60962e-19
cc_59 N_A_c_74_n N_B_XI13.X0_PGS 5.64689e-19
cc_60 N_A_c_68_n N_B_c_112_n 3.152e-19
cc_61 N_A_c_74_n N_B_c_112_n 7.5465e-19
cc_62 N_A_c_70_n N_B_c_112_n 0.00132909f
cc_63 N_A_c_70_n N_B_c_117_n 9.27569e-19
cc_64 N_Z_c_90_n N_B_c_112_n 3.31584e-19
cc_65 N_Z_c_88_n N_B_c_112_n 4.20335e-19
cc_66 N_Z_c_88_n N_B_c_117_n 0.00101313f
cc_67 N_Z_c_88_n B 0.00147455f
*
.ends
*
*
.subckt NAND2_HPNW12 A B Y VDD VSS
xgate (VSS VDD A Y B) G2_NAND2_N3
.ends
*
* File: G2_NOR2_N3.pex.netlist
* Created: Mon Feb 28 10:13:32 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_NOR2_N3_VSS 2 4 6 18 23 28 31 36 41 50 59 60 64 65 70 73 74 79 Vss
c39 74 Vss 3.75522e-19
c40 73 Vss 0.0047697f
c41 70 Vss 0.00562567f
c42 65 Vss 8.27694e-19
c43 64 Vss 0.00178035f
c44 60 Vss 6.04131e-19
c45 59 Vss 0.00565031f
c46 50 Vss 0.00520705f
c47 41 Vss 0.00279442f
c48 36 Vss 0.00113197f
c49 31 Vss 0.00124387f
c50 28 Vss 0.00807325f
c51 23 Vss 0.00817292f
c52 18 Vss 0.089128f
c53 4 Vss 0.189873f
r54 73 79 0.326018
r55 72 77 0.14525
r56 72 73 5.50157
r57 71 74 0.494161
r58 70 79 0.326018
r59 70 71 10.1279
r60 66 74 0.128424
r61 64 74 0.494161
r62 64 65 4.37625
r63 59 65 0.652036
r64 58 60 0.655813
r65 58 59 18.3386
r66 41 77 2.334
r67 36 50 1.16709
r68 36 66 2.16729
r69 31 60 1.82344
r70 28 41 1.16709
r71 23 31 1.16709
r72 16 50 0.0476429
r73 16 18 2.04225
r74 12 18 0.0685365
r75 6 28 0.123773
r76 4 12 5.1348
r77 2 23 0.123773
.ends

.subckt PM_G2_NOR2_N3_VDD 2 4 6 8 10 27 36 41 45 47 48 52 54 55 58 60 62 64 66
+ 72 78 Vss
c45 78 Vss 0.00622884f
c46 72 Vss 0.00491473f
c47 64 Vss 4.52364e-19
c48 62 Vss 0.00102348f
c49 60 Vss 6.08701e-19
c50 58 Vss 0.00198853f
c51 55 Vss 8.64913e-19
c52 54 Vss 0.00550278f
c53 52 Vss 0.0017471f
c54 49 Vss 0.0017501f
c55 48 Vss 0.00518267f
c56 47 Vss 0.00321334f
c57 45 Vss 0.0127334f
c58 41 Vss 0.00818763f
c59 37 Vss 0.129193f
c60 36 Vss 7.7089e-20
c61 27 Vss 0.0356247f
c62 26 Vss 0.102427f
c63 10 Vss 0.190932f
c64 8 Vss 0.189362f
c65 4 Vss 0.190692f
c66 2 Vss 0.191746f
r67 72 75 0.05
r68 62 78 1.16709
r69 60 66 0.326018
r70 60 62 2.16729
r71 58 75 1.16709
r72 56 58 2.95918
r73 54 66 0.326018
r74 54 55 10.1696
r75 50 64 0.0828784
r76 50 52 1.82344
r77 48 56 0.652036
r78 48 49 4.37625
r79 47 55 0.652036
r80 46 64 0.551426
r81 46 47 5.50157
r82 45 64 0.551426
r83 44 49 0.652036
r84 44 45 19.0888
r85 41 52 1.16709
r86 36 72 0.0238214
r87 36 37 2.26917
r88 33 36 2.26917
r89 29 78 0.0476429
r90 27 29 1.5171
r91 26 30 0.652036
r92 26 29 1.4004
r93 23 27 0.652036
r94 20 37 0.00605528
r95 17 33 0.00605528
r96 10 30 5.1348
r97 8 23 5.1348
r98 6 41 0.123773
r99 4 17 5.1348
r100 2 20 5.1348
.ends

.subckt PM_G2_NOR2_N3_B 2 4 10 13 18 21 26 31 Vss
c20 31 Vss 0.0033745f
c21 26 Vss 0.00378619f
c22 18 Vss 0.00118409f
c23 13 Vss 0.166574f
c24 10 Vss 7.77222e-20
c25 2 Vss 0.16675f
r26 23 31 1.16709
r27 21 23 2.37568
r28 18 26 1.16709
r29 18 21 2.45904
r30 13 31 0.50025
r31 10 26 0.50025
r32 4 13 4.37625
r33 2 10 4.37625
.ends

.subckt PM_G2_NOR2_N3_Z 2 4 6 18 22 25 28 Vss
c24 25 Vss 0.00353787f
c25 22 Vss 0.0056593f
c26 18 Vss 0.00813452f
c27 6 Vss 0.00143493f
r28 28 30 6.16843
r29 25 28 6.66857
r30 22 30 1.16709
r31 18 25 1.16709
r32 6 22 0.123773
r33 4 22 0.123773
r34 2 18 0.123773
.ends

.subckt PM_G2_NOR2_N3_A 2 4 10 11 14 18 21 Vss
c18 18 Vss 2.27081e-19
c19 14 Vss 0.2392f
c20 11 Vss 0.0348811f
c21 10 Vss 0.282285f
c22 2 Vss 0.269802f
r23 18 27 1.16709
r24 18 21 0.0416786
r25 14 27 0.05
r26 12 14 2.27565
r27 10 12 0.652036
r28 10 11 8.92755
r29 7 11 0.652036
r30 4 14 5.6016
r31 2 7 7.87725
.ends

.subckt G2_NOR2_N3  VSS VDD B Z A
*
* A	A
* Z	Z
* B	B
* VDD	VDD
* VSS	VSS
XI8.X0 N_Z_XI8.X0_D N_VDD_XI8.X0_PGD N_B_XI8.X0_CG N_VDD_XI8.X0_PGS
+ N_VSS_XI8.X0_S TIGFET_HPNW12
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_B_XI6.X0_CG N_A_XI6.X0_PGS N_VDD_XI6.X0_S
+ TIGFET_HPNW12
XI7.X0 N_Z_XI7.X0_D N_VDD_XI7.X0_PGD N_A_XI7.X0_CG N_VDD_XI7.X0_PGS
+ N_VSS_XI7.X0_S TIGFET_HPNW12
*
x_PM_G2_NOR2_N3_VSS N_VSS_XI8.X0_S N_VSS_XI6.X0_PGD N_VSS_XI7.X0_S N_VSS_c_2_p
+ N_VSS_c_8_p N_VSS_c_31_p N_VSS_c_3_p N_VSS_c_6_p N_VSS_c_32_p N_VSS_c_13_p
+ N_VSS_c_4_p N_VSS_c_5_p N_VSS_c_14_p N_VSS_c_17_p N_VSS_c_15_p N_VSS_c_20_p
+ N_VSS_c_16_p VSS Vss PM_G2_NOR2_N3_VSS
x_PM_G2_NOR2_N3_VDD N_VDD_XI8.X0_PGD N_VDD_XI8.X0_PGS N_VDD_XI6.X0_S
+ N_VDD_XI7.X0_PGD N_VDD_XI7.X0_PGS N_VDD_c_41_n N_VDD_c_63_p N_VDD_c_70_p
+ N_VDD_c_42_n N_VDD_c_45_n N_VDD_c_47_n N_VDD_c_49_n N_VDD_c_50_n N_VDD_c_56_n
+ N_VDD_c_65_p N_VDD_c_57_n N_VDD_c_58_n N_VDD_c_60_n VDD N_VDD_c_66_p
+ N_VDD_c_61_n Vss PM_G2_NOR2_N3_VDD
x_PM_G2_NOR2_N3_B N_B_XI8.X0_CG N_B_XI6.X0_CG N_B_c_90_n N_B_c_100_p N_B_c_85_n
+ B N_B_c_94_n N_B_c_88_n Vss PM_G2_NOR2_N3_B
x_PM_G2_NOR2_N3_Z N_Z_XI8.X0_D N_Z_XI6.X0_D N_Z_XI7.X0_D N_Z_c_105_n N_Z_c_107_n
+ N_Z_c_109_n Z Vss PM_G2_NOR2_N3_Z
x_PM_G2_NOR2_N3_A N_A_XI6.X0_PGS N_A_XI7.X0_CG N_A_c_129_n N_A_c_132_n
+ N_A_c_134_n N_A_c_136_n A Vss PM_G2_NOR2_N3_A
cc_1 N_VSS_XI6.X0_PGD N_VDD_XI7.X0_PGD 0.00209072f
cc_2 N_VSS_c_2_p N_VDD_c_41_n 0.00209072f
cc_3 N_VSS_c_3_p N_VDD_c_42_n 0.00187494f
cc_4 N_VSS_c_4_p N_VDD_c_42_n 0.00752502f
cc_5 N_VSS_c_5_p N_VDD_c_42_n 0.00189882f
cc_6 N_VSS_c_6_p N_VDD_c_45_n 4.76491e-19
cc_7 N_VSS_c_4_p N_VDD_c_45_n 0.00426824f
cc_8 N_VSS_c_8_p N_VDD_c_47_n 2.3316e-19
cc_9 N_VSS_c_3_p N_VDD_c_47_n 7.26139e-19
cc_10 N_VSS_c_3_p N_VDD_c_49_n 4.01154e-19
cc_11 N_VSS_c_2_p N_VDD_c_50_n 3.71132e-19
cc_12 N_VSS_c_6_p N_VDD_c_50_n 0.00141228f
cc_13 N_VSS_c_13_p N_VDD_c_50_n 0.00114511f
cc_14 N_VSS_c_14_p N_VDD_c_50_n 0.00352847f
cc_15 N_VSS_c_15_p N_VDD_c_50_n 0.00446295f
cc_16 N_VSS_c_16_p N_VDD_c_50_n 7.74609e-19
cc_17 N_VSS_c_17_p N_VDD_c_56_n 0.00106582f
cc_18 N_VSS_c_15_p N_VDD_c_57_n 0.00151536f
cc_19 N_VSS_c_6_p N_VDD_c_58_n 0.00109227f
cc_20 N_VSS_c_20_p N_VDD_c_58_n 3.86251e-19
cc_21 N_VSS_c_4_p N_VDD_c_60_n 0.00116512f
cc_22 N_VSS_c_6_p N_VDD_c_61_n 3.44698e-19
cc_23 N_VSS_c_13_p N_VDD_c_61_n 6.36088e-19
cc_24 N_VSS_c_6_p N_B_c_85_n 2.00737e-19
cc_25 N_VSS_c_13_p N_B_c_85_n 2.34295e-19
cc_26 N_VSS_c_4_p N_B_c_85_n 0.0014669f
cc_27 N_VSS_c_6_p N_B_c_88_n 2.15082e-19
cc_28 N_VSS_c_13_p N_B_c_88_n 5.20396e-19
cc_29 N_VSS_c_8_p N_Z_c_105_n 3.43419e-19
cc_30 N_VSS_c_3_p N_Z_c_105_n 3.48267e-19
cc_31 N_VSS_c_31_p N_Z_c_107_n 3.43419e-19
cc_32 N_VSS_c_32_p N_Z_c_107_n 3.48267e-19
cc_33 N_VSS_c_8_p N_Z_c_109_n 3.48267e-19
cc_34 N_VSS_c_31_p N_Z_c_109_n 3.48267e-19
cc_35 N_VSS_c_3_p N_Z_c_109_n 8.54909e-19
cc_36 N_VSS_c_32_p N_Z_c_109_n 5.71987e-19
cc_37 N_VSS_c_4_p N_Z_c_109_n 0.00105386f
cc_38 N_VSS_c_15_p N_Z_c_109_n 2.24858e-19
cc_39 N_VSS_XI6.X0_PGD N_A_c_129_n 7.89465e-19
cc_40 N_VDD_c_63_p N_B_c_90_n 4.99294e-19
cc_41 N_VDD_c_42_n N_B_c_85_n 0.0026351f
cc_42 N_VDD_c_65_p N_B_c_85_n 3.50338e-19
cc_43 N_VDD_c_66_p N_B_c_85_n 2.36346e-19
cc_44 N_VDD_c_42_n N_B_c_94_n 5.07158e-19
cc_45 N_VDD_c_65_p N_B_c_94_n 2.30903e-19
cc_46 N_VDD_c_42_n N_B_c_88_n 3.66936e-19
cc_47 N_VDD_c_70_p N_Z_c_107_n 3.43419e-19
cc_48 N_VDD_c_49_n N_Z_c_107_n 3.72199e-19
cc_49 N_VDD_c_50_n N_Z_c_107_n 2.74986e-19
cc_50 N_VDD_c_70_p N_Z_c_109_n 3.48267e-19
cc_51 N_VDD_c_42_n N_Z_c_109_n 0.00130587f
cc_52 N_VDD_c_49_n N_Z_c_109_n 7.92786e-19
cc_53 N_VDD_c_50_n N_Z_c_109_n 3.84599e-19
cc_54 N_VDD_XI8.X0_PGD N_A_c_129_n 5.98669e-19
cc_55 N_VDD_XI7.X0_PGD N_A_c_129_n 2.07763e-19
cc_56 N_VDD_XI8.X0_PGS N_A_c_132_n 8.07534e-19
cc_57 N_VDD_c_42_n N_A_c_132_n 5.64288e-19
cc_58 N_VDD_c_58_n N_A_c_134_n 2.30699e-19
cc_59 N_VDD_c_61_n N_A_c_134_n 5.11881e-19
cc_60 N_VDD_c_58_n N_A_c_136_n 2.87155e-19
cc_61 N_VDD_c_61_n N_A_c_136_n 2.16965e-19
cc_62 N_B_c_85_n N_Z_c_109_n 0.00740143f
cc_63 N_B_c_94_n N_Z_c_109_n 0.0010409f
cc_64 N_B_c_88_n N_Z_c_109_n 9.58642e-19
cc_65 N_B_c_100_p N_A_XI6.X0_PGS 4.87172e-19
cc_66 N_B_c_88_n N_A_XI6.X0_PGS 0.00109812f
cc_67 N_B_c_94_n N_A_c_129_n 0.00222679f
cc_68 N_B_c_88_n N_A_c_129_n 4.51405e-19
cc_69 N_B_c_88_n N_A_c_134_n 8.88364e-19
cc_70 N_Z_c_107_n N_A_c_129_n 4.45349e-19
cc_71 N_Z_c_109_n N_A_c_129_n 9.69188e-19
cc_72 N_Z_c_109_n N_A_c_134_n 0.00114087f
cc_73 N_Z_c_109_n N_A_c_136_n 0.00155484f
*
.ends
*
*
.subckt NOR2_HPNW12 A B Y VDD VSS
xgate (VSS VDD B Y A) G2_NOR2_N3
.ends
*
* File: G2_OAI21_N3.pex.netlist
* Created: Wed Mar  2 11:39:40 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G2_OAI21_N3_VSS 2 4 6 8 10 22 29 37 42 45 50 55 64 73 74 78 84 86 91
+ 94 Vss
c48 92 Vss 5.73928e-19
c49 91 Vss 0.00930467f
c50 86 Vss 0.00178323f
c51 84 Vss 0.00287693f
c52 79 Vss 0.00137325f
c53 78 Vss 0.00727688f
c54 74 Vss 6.08576e-19
c55 73 Vss 0.00762928f
c56 64 Vss 0.00685524f
c57 55 Vss 2.01979e-19
c58 50 Vss 0.00208662f
c59 45 Vss 0.00137663f
c60 42 Vss 0.00818763f
c61 37 Vss 0.00963114f
c62 33 Vss 0.0307825f
c63 29 Vss 5.22622e-20
c64 26 Vss 0.101261f
c65 22 Vss 0.0345879f
c66 21 Vss 0.0712517f
c67 10 Vss 0.191158f
c68 8 Vss 0.19018f
c69 4 Vss 0.189789f
r70 91 94 0.326018
r71 90 91 18.8387
r72 86 90 0.655813
r73 85 92 0.494161
r74 84 94 0.326018
r75 84 85 4.33457
r76 80 92 0.128424
r77 78 92 0.494161
r78 78 79 10.1696
r79 73 79 0.652036
r80 72 74 0.655813
r81 72 73 18.8387
r82 55 86 1.82344
r83 50 64 1.16709
r84 50 80 2.16729
r85 45 74 1.82344
r86 42 55 1.16709
r87 37 45 1.16709
r88 29 64 0.238214
r89 27 33 0.494161
r90 27 29 1.5171
r91 26 30 0.652036
r92 26 29 1.4004
r93 23 33 0.128424
r94 21 33 0.494161
r95 21 22 2.8008
r96 18 22 0.652036
r97 10 30 5.1348
r98 8 23 5.1348
r99 6 42 0.123773
r100 4 18 5.1348
r101 2 37 0.123773
.ends

.subckt PM_G2_OAI21_N3_VDD 2 4 6 8 30 35 38 39 41 43 49 51 56 59 65 Vss
c48 65 Vss 0.00671256f
c49 57 Vss 5.35171e-19
c50 56 Vss 0.0125966f
c51 55 Vss 0.0017875f
c52 51 Vss 0.00240793f
c53 49 Vss 0.00382188f
c54 47 Vss 0.00183797f
c55 43 Vss 0.00172744f
c56 41 Vss 8.2329e-19
c57 40 Vss 0.0017875f
c58 39 Vss 0.00981811f
c59 38 Vss 0.0129397f
c60 35 Vss 0.00815963f
c61 30 Vss 0.0082356f
c62 25 Vss 0.0855608f
c63 19 Vss 0.034095f
c64 18 Vss 0.0688526f
c65 6 Vss 0.192138f
c66 2 Vss 0.192543f
r67 55 59 0.326018
r68 55 56 18.8804
r69 51 56 0.655813
r70 51 53 1.82344
r71 50 57 0.494161
r72 49 59 0.326018
r73 49 50 4.37625
r74 47 65 1.16709
r75 45 57 0.128424
r76 45 47 2.20896
r77 41 43 1.82344
r78 39 57 0.494161
r79 39 40 10.1279
r80 38 41 0.655813
r81 37 40 0.652036
r82 37 38 18.8804
r83 35 53 1.16709
r84 30 43 1.16709
r85 25 65 0.238214
r86 23 25 2.04225
r87 20 23 0.0685365
r88 18 23 0.5835
r89 18 19 2.8008
r90 15 19 0.652036
r91 8 35 0.123773
r92 6 20 5.1348
r93 4 30 0.123773
r94 2 15 5.1348
.ends

.subckt PM_G2_OAI21_N3_B 2 4 13 18 21 26 31 Vss
c19 31 Vss 0.00415668f
c20 26 Vss 0.0032846f
c21 18 Vss 9.6577e-19
c22 13 Vss 0.167996f
c23 2 Vss 0.166757f
r24 23 31 1.16709
r25 21 23 1.66714
r26 18 26 1.16709
r27 18 21 3.16757
r28 13 31 0.476429
r29 10 26 0.50025
r30 4 13 4.4346
r31 2 10 4.37625
.ends

.subckt PM_G2_OAI21_N3_A 2 4 13 18 21 26 31 36 44 46 Vss
c38 46 Vss 1.44014e-19
c39 36 Vss 0.00294987f
c40 31 Vss 0.00806931f
c41 26 Vss 0.0038514f
c42 21 Vss 0.00314266f
c43 18 Vss 0.0859029f
c44 13 Vss 4.64808e-20
c45 4 Vss 0.166608f
c46 2 Vss 0.193159f
r47 40 46 0.655813
r48 26 36 1.16709
r49 26 46 4.52212
r50 21 31 1.16709
r51 21 44 0.0833571
r52 21 40 12.6703
r53 18 31 0.238214
r54 15 18 1.92555
r55 13 36 0.50025
r56 7 15 0.0685365
r57 4 13 4.37625
r58 2 7 5.1348
.ends

.subckt PM_G2_OAI21_N3_Z 2 4 6 8 23 27 30 33 Vss
c33 30 Vss 0.0016158f
c34 27 Vss 0.00640524f
c35 23 Vss 0.00630974f
c36 8 Vss 0.00143493f
c37 6 Vss 0.00143493f
r38 33 35 7.54382
r39 30 33 5.29318
r40 27 35 1.16709
r41 23 30 1.16709
r42 8 27 0.123773
r43 6 23 0.123773
r44 4 27 0.123773
r45 2 23 0.123773
.ends

.subckt PM_G2_OAI21_N3_C 2 4 6 13 14 17 24 27 Vss
c28 27 Vss 7.80628e-19
c29 24 Vss 0.0813012f
c30 17 Vss 0.25734f
c31 14 Vss 0.0348849f
c32 13 Vss 0.247183f
c33 4 Vss 0.29011f
c34 2 Vss 0.290309f
r35 27 30 0.0833571
r36 23 24 2.04225
r37 20 24 0.0685365
r38 17 30 1.16709
r39 15 23 0.0685365
r40 15 17 2.8008
r41 13 23 0.5835
r42 13 14 8.92755
r43 10 14 0.652036
r44 6 17 5.6016
r45 4 20 8.4024
r46 2 10 8.4024
.ends

.subckt G2_OAI21_N3  VSS VDD B A Z C
*
* C	C
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI7.X0 N_Z_XI7.X0_D N_VDD_XI7.X0_PGD N_B_XI7.X0_CG N_C_XI7.X0_PGS N_VSS_XI7.X0_S
+ TIGFET_HPNW12
XI5.X0 N_Z_XI5.X0_D N_VSS_XI5.X0_PGD N_B_XI5.X0_CG N_A_XI5.X0_PGS N_VDD_XI5.X0_S
+ TIGFET_HPNW12
XI8.X0 N_Z_XI8.X0_D N_VDD_XI8.X0_PGD N_A_XI8.X0_CG N_C_XI8.X0_PGS N_VSS_XI8.X0_S
+ TIGFET_HPNW12
XI6.X0 N_Z_XI6.X0_D N_VSS_XI6.X0_PGD N_C_XI6.X0_CG N_VSS_XI6.X0_PGS
+ N_VDD_XI6.X0_S TIGFET_HPNW12
*
x_PM_G2_OAI21_N3_VSS N_VSS_XI7.X0_S N_VSS_XI5.X0_PGD N_VSS_XI8.X0_S
+ N_VSS_XI6.X0_PGD N_VSS_XI6.X0_PGS N_VSS_c_30_p N_VSS_c_46_p N_VSS_c_1_p
+ N_VSS_c_10_p N_VSS_c_2_p N_VSS_c_22_p N_VSS_c_11_p N_VSS_c_23_p N_VSS_c_3_p
+ N_VSS_c_4_p N_VSS_c_9_p N_VSS_c_13_p N_VSS_c_12_p N_VSS_c_15_p VSS Vss
+ PM_G2_OAI21_N3_VSS
x_PM_G2_OAI21_N3_VDD N_VDD_XI7.X0_PGD N_VDD_XI5.X0_S N_VDD_XI8.X0_PGD
+ N_VDD_XI6.X0_S N_VDD_c_80_p N_VDD_c_81_p N_VDD_c_49_n N_VDD_c_53_n
+ N_VDD_c_55_n N_VDD_c_56_n N_VDD_c_58_n N_VDD_c_61_n N_VDD_c_64_n VDD
+ N_VDD_c_71_p Vss PM_G2_OAI21_N3_VDD
x_PM_G2_OAI21_N3_B N_B_XI7.X0_CG N_B_XI5.X0_CG N_B_c_103_p N_B_c_97_n B
+ N_B_c_99_n N_B_c_100_n Vss PM_G2_OAI21_N3_B
x_PM_G2_OAI21_N3_A N_A_XI5.X0_PGS N_A_XI8.X0_CG N_A_c_130_n N_A_c_137_n
+ N_A_c_117_n N_A_c_122_n N_A_c_124_n N_A_c_134_n A N_A_c_128_n Vss
+ PM_G2_OAI21_N3_A
x_PM_G2_OAI21_N3_Z N_Z_XI7.X0_D N_Z_XI5.X0_D N_Z_XI8.X0_D N_Z_XI6.X0_D
+ N_Z_c_154_n N_Z_c_165_n N_Z_c_158_n Z Vss PM_G2_OAI21_N3_Z
x_PM_G2_OAI21_N3_C N_C_XI7.X0_PGS N_C_XI8.X0_PGS N_C_XI6.X0_CG N_C_c_187_n
+ N_C_c_206_n N_C_c_189_n N_C_c_191_n C Vss PM_G2_OAI21_N3_C
cc_1 N_VSS_c_1_p N_VDD_c_49_n 9.5668e-19
cc_2 N_VSS_c_2_p N_VDD_c_49_n 0.00165395f
cc_3 N_VSS_c_3_p N_VDD_c_49_n 0.00820308f
cc_4 N_VSS_c_4_p N_VDD_c_49_n 0.00189979f
cc_5 N_VSS_c_1_p N_VDD_c_53_n 2.43883e-19
cc_6 N_VSS_c_2_p N_VDD_c_53_n 7.51487e-19
cc_7 N_VSS_c_3_p N_VDD_c_55_n 0.00170274f
cc_8 N_VSS_c_2_p N_VDD_c_56_n 4.01889e-19
cc_9 N_VSS_c_9_p N_VDD_c_56_n 4.74109e-19
cc_10 N_VSS_c_10_p N_VDD_c_58_n 2.43883e-19
cc_11 N_VSS_c_11_p N_VDD_c_58_n 3.33988e-19
cc_12 N_VSS_c_12_p N_VDD_c_58_n 4.17499e-19
cc_13 N_VSS_c_13_p N_VDD_c_61_n 4.74109e-19
cc_14 N_VSS_c_12_p N_VDD_c_61_n 4.01889e-19
cc_15 N_VSS_c_15_p N_VDD_c_61_n 0.00178085f
cc_16 N_VSS_c_10_p N_VDD_c_64_n 9.5668e-19
cc_17 N_VSS_c_11_p N_VDD_c_64_n 0.00165395f
cc_18 N_VSS_c_12_p N_VDD_c_64_n 0.00189979f
cc_19 N_VSS_c_15_p N_VDD_c_64_n 0.0087982f
cc_20 N_VSS_c_3_p N_B_c_97_n 5.69535e-19
cc_21 N_VSS_XI5.X0_PGD N_A_XI5.X0_PGS 0.00176902f
cc_22 N_VSS_c_22_p N_A_c_117_n 8.59446e-19
cc_23 N_VSS_c_23_p N_A_c_117_n 3.44698e-19
cc_24 N_VSS_c_3_p N_A_c_117_n 0.00485346f
cc_25 N_VSS_c_9_p N_A_c_117_n 0.00211426f
cc_26 N_VSS_c_15_p N_A_c_117_n 0.00226606f
cc_27 N_VSS_c_9_p N_A_c_122_n 6.38907e-19
cc_28 N_VSS_c_15_p N_A_c_122_n 7.9739e-19
cc_29 N_VSS_XI5.X0_PGD N_A_c_124_n 3.11814e-19
cc_30 N_VSS_c_30_p N_A_c_124_n 0.00322564f
cc_31 N_VSS_c_22_p N_A_c_124_n 3.44698e-19
cc_32 N_VSS_c_23_p N_A_c_124_n 6.61253e-19
cc_33 N_VSS_c_3_p N_A_c_128_n 0.00309992f
cc_34 N_VSS_c_1_p N_Z_c_154_n 3.43419e-19
cc_35 N_VSS_c_10_p N_Z_c_154_n 3.43419e-19
cc_36 N_VSS_c_2_p N_Z_c_154_n 3.48267e-19
cc_37 N_VSS_c_11_p N_Z_c_154_n 3.48267e-19
cc_38 N_VSS_c_1_p N_Z_c_158_n 3.48267e-19
cc_39 N_VSS_c_10_p N_Z_c_158_n 3.48267e-19
cc_40 N_VSS_c_2_p N_Z_c_158_n 5.71987e-19
cc_41 N_VSS_c_11_p N_Z_c_158_n 5.71987e-19
cc_42 N_VSS_c_9_p N_Z_c_158_n 3.21537e-19
cc_43 N_VSS_c_15_p N_Z_c_158_n 8.14216e-19
cc_44 N_VSS_XI5.X0_PGD N_C_c_187_n 6.83817e-19
cc_45 N_VSS_XI6.X0_PGD N_C_c_187_n 6.83817e-19
cc_46 N_VSS_c_46_p N_C_c_189_n 2.53848e-19
cc_47 N_VSS_c_23_p N_C_c_189_n 0.00232974f
cc_48 N_VSS_XI6.X0_PGS N_C_c_191_n 8.42974e-19
cc_49 N_VDD_c_49_n N_B_c_97_n 0.00231792f
cc_50 N_VDD_c_49_n N_B_c_99_n 3.66936e-19
cc_51 N_VDD_c_49_n N_B_c_100_n 4.8547e-19
cc_52 N_VDD_c_71_p N_A_XI8.X0_CG 0.00266603f
cc_53 N_VDD_c_71_p N_A_c_130_n 5.2106e-19
cc_54 N_VDD_c_53_n N_A_c_122_n 6.20865e-19
cc_55 N_VDD_c_64_n N_A_c_122_n 6.23587e-19
cc_56 N_VDD_c_71_p N_A_c_122_n 2.23358e-19
cc_57 N_VDD_c_64_n N_A_c_134_n 3.66936e-19
cc_58 N_VDD_c_71_p N_A_c_134_n 3.65437e-19
cc_59 N_VDD_c_49_n N_A_c_128_n 6.11072e-19
cc_60 N_VDD_c_53_n N_Z_c_154_n 2.43883e-19
cc_61 N_VDD_c_80_p N_Z_c_165_n 3.43419e-19
cc_62 N_VDD_c_81_p N_Z_c_165_n 3.43419e-19
cc_63 N_VDD_c_56_n N_Z_c_165_n 3.72199e-19
cc_64 N_VDD_c_61_n N_Z_c_165_n 3.72199e-19
cc_65 N_VDD_c_80_p N_Z_c_158_n 3.48267e-19
cc_66 N_VDD_c_81_p N_Z_c_158_n 3.48267e-19
cc_67 N_VDD_c_49_n N_Z_c_158_n 0.00116129f
cc_68 N_VDD_c_53_n N_Z_c_158_n 5.05821e-19
cc_69 N_VDD_c_56_n N_Z_c_158_n 5.09542e-19
cc_70 N_VDD_c_61_n N_Z_c_158_n 7.72285e-19
cc_71 N_VDD_c_64_n N_Z_c_158_n 0.00182594f
cc_72 N_VDD_c_49_n N_C_XI7.X0_PGS 6.13097e-19
cc_73 N_VDD_c_64_n N_C_XI8.X0_PGS 6.32546e-19
cc_74 N_VDD_XI7.X0_PGD N_C_c_187_n 6.83817e-19
cc_75 N_VDD_XI8.X0_PGD N_C_c_187_n 6.83817e-19
cc_76 N_VDD_c_64_n N_C_c_189_n 5.92666e-19
cc_77 N_VDD_c_64_n C 5.04211e-19
cc_78 N_B_c_100_n N_A_c_137_n 2.60115e-19
cc_79 N_B_c_97_n N_A_c_117_n 0.00265561f
cc_80 N_B_c_103_p N_A_c_124_n 0.00262973f
cc_81 N_B_c_97_n N_A_c_124_n 2.40146e-19
cc_82 N_B_c_100_n N_A_c_124_n 3.65437e-19
cc_83 N_B_c_99_n N_A_c_134_n 8.86454e-19
cc_84 N_B_c_97_n N_A_c_128_n 7.49556e-19
cc_85 N_B_c_97_n N_Z_c_158_n 0.00671f
cc_86 N_B_c_99_n N_Z_c_158_n 9.58174e-19
cc_87 N_B_c_100_n N_Z_c_158_n 0.00101748f
cc_88 N_B_XI7.X0_CG N_C_XI7.X0_PGS 4.87172e-19
cc_89 N_B_c_99_n N_C_XI7.X0_PGS 0.001089f
cc_90 N_B_c_99_n N_C_c_187_n 6.02551e-19
cc_91 N_B_c_100_n N_C_c_187_n 0.00149356f
cc_92 N_B_c_100_n N_C_c_189_n 9.54365e-19
cc_93 N_A_c_117_n N_Z_c_158_n 0.00195546f
cc_94 N_A_c_122_n N_Z_c_158_n 0.00358051f
cc_95 N_A_c_134_n N_Z_c_158_n 9.53427e-19
cc_96 N_A_XI8.X0_CG N_C_XI8.X0_PGS 4.87172e-19
cc_97 N_A_c_134_n N_C_XI8.X0_PGS 0.001089f
cc_98 N_A_c_134_n N_C_c_187_n 0.00157146f
cc_99 N_A_XI5.X0_PGS N_C_c_206_n 8.42974e-19
cc_100 N_A_c_122_n N_C_c_189_n 5.38228e-19
cc_101 N_A_c_134_n N_C_c_189_n 0.00222154f
cc_102 N_A_c_122_n C 8.18489e-19
cc_103 N_Z_c_154_n N_C_c_187_n 3.5202e-19
cc_104 N_Z_c_165_n N_C_c_187_n 3.5202e-19
cc_105 N_Z_c_158_n N_C_c_187_n 3.56555e-19
cc_106 N_Z_c_158_n N_C_c_189_n 0.00101565f
cc_107 N_Z_c_158_n C 0.00141616f
*
.ends
*
*
.subckt OAI21_HPNW12 A0 A1 B0 Y VDD VSS
xgate (VSS VDD A1 A0 Y B0) G2_OAI21_N3
.ends
*
* File: G3_OR2_N3.pex.netlist
* Created: Tue Mar  1 12:18:46 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G3_OR2_N3_VSS 2 4 6 8 10 12 28 29 38 44 49 52 57 62 67 76 85 90 91 95
+ 96 101 107 114 115 116 Vss
c71 116 Vss 3.91906e-19
c72 115 Vss 3.75522e-19
c73 107 Vss 0.00372185f
c74 101 Vss 0.00290457f
c75 96 Vss 8.35017e-19
c76 95 Vss 0.00178035f
c77 91 Vss 6.20207e-19
c78 90 Vss 0.00579798f
c79 85 Vss 0.0039758f
c80 76 Vss 0.0050462f
c81 67 Vss 5.89061e-19
c82 62 Vss 8.97934e-19
c83 57 Vss 0.00103095f
c84 52 Vss 0.00124124f
c85 49 Vss 0.00687623f
c86 44 Vss 0.00812495f
c87 38 Vss 0.0895788f
c88 29 Vss 0.0349332f
c89 28 Vss 0.0997249f
c90 12 Vss 0.190073f
c91 10 Vss 0.189045f
c92 8 Vss 0.00143493f
c93 4 Vss 0.189407f
r94 109 114 0.458464
r95 108 116 0.494161
r96 107 109 0.652036
r97 107 108 7.46046
r98 103 116 0.128424
r99 102 115 0.494161
r100 101 116 0.494161
r101 101 102 7.46046
r102 97 115 0.128424
r103 95 115 0.494161
r104 95 96 4.37625
r105 90 96 0.652036
r106 89 91 0.655813
r107 89 90 18.3386
r108 67 85 1.16709
r109 67 114 1.70882
r110 62 103 6.16843
r111 57 76 1.16709
r112 57 97 2.16729
r113 52 91 1.82344
r114 49 62 1.16709
r115 44 52 1.16709
r116 36 76 0.0476429
r117 36 38 2.04225
r118 31 85 0.0476429
r119 29 31 1.45875
r120 28 32 0.652036
r121 28 31 1.45875
r122 25 29 0.652036
r123 22 38 0.0685365
r124 12 32 5.1348
r125 10 25 5.1348
r126 8 49 0.123773
r127 6 49 0.123773
r128 4 22 5.1348
r129 2 44 0.123773
.ends

.subckt PM_G3_OR2_N3_VDD 2 4 6 8 10 12 14 16 37 46 56 62 67 70 72 73 77 79 80 83
+ 87 89 93 95 97 102 103 104 105 107 113 119 124 Vss
c78 124 Vss 0.00450608f
c79 119 Vss 0.00587228f
c80 113 Vss 0.00493107f
c81 105 Vss 2.39889e-19
c82 104 Vss 2.39889e-19
c83 103 Vss 4.52364e-19
c84 102 Vss 0.00430335f
c85 101 Vss 0.00170674f
c86 97 Vss 0.00160078f
c87 95 Vss 0.00854117f
c88 93 Vss 7.28478e-19
c89 89 Vss 0.00205766f
c90 87 Vss 4.80319e-19
c91 83 Vss 0.00133062f
c92 80 Vss 8.68835e-19
c93 79 Vss 0.00561215f
c94 77 Vss 0.0017471f
c95 74 Vss 0.00174847f
c96 73 Vss 0.00498635f
c97 72 Vss 0.00313638f
c98 70 Vss 0.0119561f
c99 67 Vss 0.0100342f
c100 62 Vss 0.00818522f
c101 57 Vss 0.129193f
c102 56 Vss 7.73513e-20
c103 47 Vss 0.035874f
c104 46 Vss 0.101312f
c105 37 Vss 0.0356247f
c106 36 Vss 0.101564f
c107 14 Vss 0.189069f
c108 12 Vss 0.189513f
c109 10 Vss 0.189312f
c110 8 Vss 0.189362f
c111 4 Vss 0.191197f
c112 2 Vss 0.192293f
r113 113 116 0.05
r114 101 107 0.349767
r115 101 102 5.50157
r116 97 107 0.306046
r117 97 99 1.82344
r118 96 105 0.494161
r119 95 102 0.652036
r120 95 96 10.1279
r121 93 124 1.16709
r122 91 105 0.128424
r123 91 93 2.16729
r124 90 104 0.494161
r125 89 105 0.494161
r126 89 90 4.54296
r127 87 119 1.16709
r128 85 104 0.128424
r129 85 87 2.16729
r130 83 116 1.16709
r131 81 83 2.16729
r132 79 104 0.494161
r133 79 80 10.1696
r134 75 103 0.0828784
r135 75 77 1.82344
r136 73 81 0.652036
r137 73 74 4.37625
r138 72 80 0.652036
r139 71 103 0.551426
r140 71 72 5.50157
r141 70 103 0.551426
r142 69 74 0.652036
r143 69 70 18.2969
r144 67 99 1.16709
r145 62 77 1.16709
r146 56 113 0.0238214
r147 56 57 2.26917
r148 53 56 2.26917
r149 49 124 0.0476429
r150 47 49 1.45875
r151 46 50 0.652036
r152 46 49 1.45875
r153 43 47 0.652036
r154 39 119 0.0476429
r155 37 39 1.5171
r156 36 40 0.652036
r157 36 39 1.4004
r158 33 37 0.652036
r159 30 57 0.00605528
r160 27 53 0.00605528
r161 16 67 0.123773
r162 14 43 5.1348
r163 12 50 5.1348
r164 10 40 5.1348
r165 8 33 5.1348
r166 6 62 0.123773
r167 4 27 5.1348
r168 2 30 5.1348
.ends

.subckt PM_G3_OR2_N3_B 2 4 10 13 18 21 26 31 Vss
c19 31 Vss 0.00192399f
c20 26 Vss 0.00378619f
c21 18 Vss 0.00125219f
c22 13 Vss 0.166574f
c23 10 Vss 7.84101e-20
c24 2 Vss 0.16675f
r25 23 31 1.16709
r26 21 23 2.29232
r27 18 26 1.16709
r28 18 21 2.54239
r29 13 31 0.50025
r30 10 26 0.50025
r31 4 13 4.37625
r32 2 10 4.37625
.ends

.subckt PM_G3_OR2_N3_NET21 2 4 6 8 10 24 27 38 42 45 53 66 70 Vss
c35 70 Vss 0.00748471f
c36 66 Vss 0.00592889f
c37 53 Vss 0.0020112f
c38 45 Vss 0.00308864f
c39 42 Vss 0.00545637f
c40 38 Vss 0.00813452f
c41 27 Vss 8.95828e-20
c42 24 Vss 0.229828f
c43 21 Vss 0.18045f
c44 19 Vss 0.0247918f
c45 10 Vss 0.193588f
c46 6 Vss 0.00143493f
r47 70 74 0.652036
r48 53 66 1.16709
r49 53 74 2.16729
r50 48 70 8.04396
r51 48 50 6.75193
r52 45 48 6.08507
r53 42 50 1.16709
r54 38 45 1.16709
r55 27 66 0.0476429
r56 25 27 0.326018
r57 25 27 0.1167
r58 24 28 0.652036
r59 24 27 6.7686
r60 21 66 0.357321
r61 19 27 0.326018
r62 19 21 0.40845
r63 10 28 5.1348
r64 8 21 4.72635
r65 6 42 0.123773
r66 4 42 0.123773
r67 2 38 0.123773
.ends

.subckt PM_G3_OR2_N3_A 2 4 10 11 14 18 21 Vss
c21 18 Vss 3.08468e-19
c22 14 Vss 0.225307f
c23 11 Vss 0.0348763f
c24 10 Vss 0.278488f
c25 2 Vss 0.253009f
r26 18 27 1.16709
r27 18 21 0.0416786
r28 14 27 0.05
r29 12 14 1.6338
r30 10 12 0.652036
r31 10 11 8.92755
r32 7 11 0.652036
r33 4 14 5.6016
r34 2 7 7.2354
.ends

.subckt PM_G3_OR2_N3_Z 2 4 13 19 Vss
c12 13 Vss 0.00498872f
c13 4 Vss 0.00143493f
r14 16 19 0.0364688
r15 13 16 1.16709
r16 4 13 0.123773
r17 2 13 0.123773
.ends

.subckt G3_OR2_N3  VSS VDD B A Z
*
* Z	Z
* A	A
* B	B
* VDD	VDD
* VSS	VSS
XI12.X0 N_NET21_XI12.X0_D N_VDD_XI12.X0_PGD N_B_XI12.X0_CG N_VDD_XI12.X0_PGS
+ N_VSS_XI12.X0_S TIGFET_HPNW12
XI10.X0 N_NET21_XI10.X0_D N_VSS_XI10.X0_PGD N_B_XI10.X0_CG N_A_XI10.X0_PGS
+ N_VDD_XI10.X0_S TIGFET_HPNW12
XI11.X0 N_NET21_XI11.X0_D N_VDD_XI11.X0_PGD N_A_XI11.X0_CG N_VDD_XI11.X0_PGS
+ N_VSS_XI11.X0_S TIGFET_HPNW12
XI14.X0 N_Z_XI14.X0_D N_VDD_XI14.X0_PGD N_NET21_XI14.X0_CG N_VDD_XI14.X0_PGS
+ N_VSS_XI14.X0_S TIGFET_HPNW12
XI13.X0 N_Z_XI13.X0_D N_VSS_XI13.X0_PGD N_NET21_XI13.X0_CG N_VSS_XI13.X0_PGS
+ N_VDD_XI13.X0_S TIGFET_HPNW12
*
x_PM_G3_OR2_N3_VSS N_VSS_XI12.X0_S N_VSS_XI10.X0_PGD N_VSS_XI11.X0_S
+ N_VSS_XI14.X0_S N_VSS_XI13.X0_PGD N_VSS_XI13.X0_PGS N_VSS_c_32_p N_VSS_c_4_p
+ N_VSS_c_3_p N_VSS_c_11_p N_VSS_c_24_p N_VSS_c_5_p N_VSS_c_8_p N_VSS_c_22_p
+ N_VSS_c_30_p N_VSS_c_9_p N_VSS_c_31_p N_VSS_c_6_p N_VSS_c_7_p N_VSS_c_17_p
+ N_VSS_c_20_p N_VSS_c_18_p N_VSS_c_27_p VSS N_VSS_c_19_p N_VSS_c_28_p Vss
+ PM_G3_OR2_N3_VSS
x_PM_G3_OR2_N3_VDD N_VDD_XI12.X0_PGD N_VDD_XI12.X0_PGS N_VDD_XI10.X0_S
+ N_VDD_XI11.X0_PGD N_VDD_XI11.X0_PGS N_VDD_XI14.X0_PGD N_VDD_XI14.X0_PGS
+ N_VDD_XI13.X0_S N_VDD_c_74_n N_VDD_c_75_n N_VDD_c_119_p N_VDD_c_128_p
+ N_VDD_c_144_p N_VDD_c_76_n N_VDD_c_79_n N_VDD_c_82_n N_VDD_c_84_n N_VDD_c_85_n
+ N_VDD_c_91_n N_VDD_c_121_p N_VDD_c_92_n N_VDD_c_95_n N_VDD_c_100_n
+ N_VDD_c_103_n N_VDD_c_146_p N_VDD_c_108_n N_VDD_c_112_n N_VDD_c_113_n
+ N_VDD_c_114_n VDD N_VDD_c_122_p N_VDD_c_115_n N_VDD_c_117_n Vss
+ PM_G3_OR2_N3_VDD
x_PM_G3_OR2_N3_B N_B_XI12.X0_CG N_B_XI10.X0_CG N_B_c_155_n N_B_c_165_p
+ N_B_c_150_n B N_B_c_159_n N_B_c_153_n Vss PM_G3_OR2_N3_B
x_PM_G3_OR2_N3_NET21 N_NET21_XI12.X0_D N_NET21_XI10.X0_D N_NET21_XI11.X0_D
+ N_NET21_XI14.X0_CG N_NET21_XI13.X0_CG N_NET21_c_169_n N_NET21_c_183_n
+ N_NET21_c_170_n N_NET21_c_172_n N_NET21_c_174_n N_NET21_c_191_n
+ N_NET21_c_199_p N_NET21_c_179_n Vss PM_G3_OR2_N3_NET21
x_PM_G3_OR2_N3_A N_A_XI10.X0_PGS N_A_XI11.X0_CG N_A_c_204_n N_A_c_207_n
+ N_A_c_209_n N_A_c_211_n A Vss PM_G3_OR2_N3_A
x_PM_G3_OR2_N3_Z N_Z_XI14.X0_D N_Z_XI13.X0_D N_Z_c_225_n Z Vss PM_G3_OR2_N3_Z
cc_1 N_VSS_XI10.X0_PGD N_VDD_XI11.X0_PGD 0.00203999f
cc_2 N_VSS_XI13.X0_PGD N_VDD_XI14.X0_PGD 0.00196229f
cc_3 N_VSS_c_3_p N_VDD_c_74_n 0.00203999f
cc_4 N_VSS_c_4_p N_VDD_c_75_n 0.00196229f
cc_5 N_VSS_c_5_p N_VDD_c_76_n 0.00187494f
cc_6 N_VSS_c_6_p N_VDD_c_76_n 0.0079127f
cc_7 N_VSS_c_7_p N_VDD_c_76_n 0.00189882f
cc_8 N_VSS_c_8_p N_VDD_c_79_n 4.35319e-19
cc_9 N_VSS_c_9_p N_VDD_c_79_n 4.7255e-19
cc_10 N_VSS_c_6_p N_VDD_c_79_n 0.00412661f
cc_11 N_VSS_c_11_p N_VDD_c_82_n 2.77593e-19
cc_12 N_VSS_c_5_p N_VDD_c_82_n 8.30039e-19
cc_13 N_VSS_c_5_p N_VDD_c_84_n 4.01154e-19
cc_14 N_VSS_c_3_p N_VDD_c_85_n 3.71132e-19
cc_15 N_VSS_c_8_p N_VDD_c_85_n 0.00141228f
cc_16 N_VSS_c_9_p N_VDD_c_85_n 0.00114511f
cc_17 N_VSS_c_17_p N_VDD_c_85_n 0.00352847f
cc_18 N_VSS_c_18_p N_VDD_c_85_n 0.00442704f
cc_19 N_VSS_c_19_p N_VDD_c_85_n 7.74609e-19
cc_20 N_VSS_c_20_p N_VDD_c_91_n 0.00107113f
cc_21 N_VSS_c_8_p N_VDD_c_92_n 8.39054e-19
cc_22 N_VSS_c_22_p N_VDD_c_92_n 3.93845e-19
cc_23 N_VSS_c_9_p N_VDD_c_92_n 3.95933e-19
cc_24 N_VSS_c_24_p N_VDD_c_95_n 2.74986e-19
cc_25 N_VSS_c_22_p N_VDD_c_95_n 2.9533e-19
cc_26 N_VSS_c_18_p N_VDD_c_95_n 0.00139286f
cc_27 N_VSS_c_27_p N_VDD_c_95_n 0.0014416f
cc_28 N_VSS_c_28_p N_VDD_c_95_n 0.00111918f
cc_29 N_VSS_c_22_p N_VDD_c_100_n 3.91951e-19
cc_30 N_VSS_c_30_p N_VDD_c_100_n 8.45954e-19
cc_31 N_VSS_c_31_p N_VDD_c_100_n 3.99794e-19
cc_32 N_VSS_c_32_p N_VDD_c_103_n 4.0633e-19
cc_33 N_VSS_c_4_p N_VDD_c_103_n 3.89167e-19
cc_34 N_VSS_c_30_p N_VDD_c_103_n 0.00161703f
cc_35 N_VSS_c_31_p N_VDD_c_103_n 2.26455e-19
cc_36 N_VSS_c_27_p N_VDD_c_103_n 0.00619092f
cc_37 N_VSS_XI13.X0_PGS N_VDD_c_108_n 4.28478e-19
cc_38 N_VSS_c_22_p N_VDD_c_108_n 2.85882e-19
cc_39 N_VSS_c_30_p N_VDD_c_108_n 8.67538e-19
cc_40 N_VSS_c_31_p N_VDD_c_108_n 3.66936e-19
cc_41 N_VSS_c_6_p N_VDD_c_112_n 0.00116512f
cc_42 N_VSS_c_18_p N_VDD_c_113_n 0.00102637f
cc_43 N_VSS_c_27_p N_VDD_c_114_n 0.00103008f
cc_44 N_VSS_c_8_p N_VDD_c_115_n 3.44698e-19
cc_45 N_VSS_c_9_p N_VDD_c_115_n 6.36088e-19
cc_46 N_VSS_c_30_p N_VDD_c_117_n 3.48267e-19
cc_47 N_VSS_c_31_p N_VDD_c_117_n 6.489e-19
cc_48 N_VSS_c_8_p N_B_c_150_n 2.0198e-19
cc_49 N_VSS_c_9_p N_B_c_150_n 2.34295e-19
cc_50 N_VSS_c_6_p N_B_c_150_n 9.20502e-19
cc_51 N_VSS_c_8_p N_B_c_153_n 2.15082e-19
cc_52 N_VSS_c_9_p N_B_c_153_n 5.28949e-19
cc_53 N_VSS_XI13.X0_PGD N_NET21_c_169_n 4.31283e-19
cc_54 N_VSS_c_11_p N_NET21_c_170_n 3.43419e-19
cc_55 N_VSS_c_5_p N_NET21_c_170_n 3.48267e-19
cc_56 N_VSS_c_24_p N_NET21_c_172_n 3.43419e-19
cc_57 N_VSS_c_22_p N_NET21_c_172_n 3.48267e-19
cc_58 N_VSS_c_11_p N_NET21_c_174_n 3.48267e-19
cc_59 N_VSS_c_24_p N_NET21_c_174_n 3.48267e-19
cc_60 N_VSS_c_5_p N_NET21_c_174_n 8.54909e-19
cc_61 N_VSS_c_22_p N_NET21_c_174_n 5.71987e-19
cc_62 N_VSS_c_6_p N_NET21_c_174_n 9.99273e-19
cc_63 N_VSS_c_22_p N_NET21_c_179_n 8.10259e-19
cc_64 N_VSS_c_6_p N_NET21_c_179_n 2.03357e-19
cc_65 N_VSS_c_18_p N_NET21_c_179_n 6.96588e-19
cc_66 N_VSS_XI10.X0_PGD N_A_c_204_n 9.58706e-19
cc_67 N_VSS_c_24_p N_Z_c_225_n 3.43419e-19
cc_68 N_VSS_c_22_p N_Z_c_225_n 3.48267e-19
cc_69 N_VSS_c_24_p Z 3.48267e-19
cc_70 N_VSS_c_22_p Z 7.85754e-19
cc_71 N_VSS_c_27_p Z 2.23989e-19
cc_72 N_VDD_c_119_p N_B_c_155_n 5.04908e-19
cc_73 N_VDD_c_76_n N_B_c_150_n 0.00268701f
cc_74 N_VDD_c_121_p N_B_c_150_n 3.49578e-19
cc_75 N_VDD_c_122_p N_B_c_150_n 2.36346e-19
cc_76 N_VDD_c_76_n N_B_c_159_n 5.07158e-19
cc_77 N_VDD_c_121_p N_B_c_159_n 2.30699e-19
cc_78 N_VDD_c_76_n N_B_c_153_n 3.66936e-19
cc_79 N_VDD_XI14.X0_PGD N_NET21_c_169_n 4.31283e-19
cc_80 N_VDD_c_117_n N_NET21_c_183_n 5.33384e-19
cc_81 N_VDD_c_128_p N_NET21_c_172_n 3.43419e-19
cc_82 N_VDD_c_84_n N_NET21_c_172_n 3.72199e-19
cc_83 N_VDD_c_85_n N_NET21_c_172_n 2.74986e-19
cc_84 N_VDD_c_128_p N_NET21_c_174_n 3.48267e-19
cc_85 N_VDD_c_76_n N_NET21_c_174_n 0.00123401f
cc_86 N_VDD_c_84_n N_NET21_c_174_n 7.92786e-19
cc_87 N_VDD_c_85_n N_NET21_c_174_n 3.84599e-19
cc_88 N_VDD_c_117_n N_NET21_c_191_n 2.15082e-19
cc_89 N_VDD_XI12.X0_PGD N_A_c_204_n 5.14897e-19
cc_90 N_VDD_XI11.X0_PGD N_A_c_204_n 2.52296e-19
cc_91 N_VDD_XI12.X0_PGS N_A_c_207_n 6.93093e-19
cc_92 N_VDD_c_76_n N_A_c_207_n 5.08654e-19
cc_93 N_VDD_c_92_n N_A_c_209_n 2.30699e-19
cc_94 N_VDD_c_115_n N_A_c_209_n 5.05291e-19
cc_95 N_VDD_c_92_n N_A_c_211_n 2.64342e-19
cc_96 N_VDD_c_115_n N_A_c_211_n 2.15082e-19
cc_97 N_VDD_c_144_p N_Z_c_225_n 3.43419e-19
cc_98 N_VDD_c_103_n N_Z_c_225_n 2.74986e-19
cc_99 N_VDD_c_146_p N_Z_c_225_n 3.72199e-19
cc_100 N_VDD_c_144_p Z 3.48267e-19
cc_101 N_VDD_c_103_n Z 3.66281e-19
cc_102 N_VDD_c_146_p Z 7.4527e-19
cc_103 N_B_c_150_n N_NET21_c_174_n 0.00754318f
cc_104 N_B_c_159_n N_NET21_c_174_n 0.0010409f
cc_105 N_B_c_153_n N_NET21_c_174_n 9.33005e-19
cc_106 N_B_c_165_p N_A_XI10.X0_PGS 4.87172e-19
cc_107 N_B_c_153_n N_A_XI10.X0_PGS 7.86826e-19
cc_108 N_B_c_159_n N_A_c_204_n 0.00191474f
cc_109 N_B_c_153_n N_A_c_209_n 7.50183e-19
cc_110 N_NET21_c_172_n N_A_c_204_n 4.90018e-19
cc_111 N_NET21_c_174_n N_A_c_204_n 8.56417e-19
cc_112 N_NET21_c_174_n N_A_c_209_n 0.00108943f
cc_113 N_NET21_c_191_n N_A_c_209_n 3.48267e-19
cc_114 N_NET21_c_199_p N_A_c_209_n 0.00171208f
cc_115 N_NET21_c_174_n N_A_c_211_n 0.00142917f
cc_116 N_NET21_c_191_n N_A_c_211_n 4.28721e-19
cc_117 N_NET21_c_179_n N_A_c_211_n 3.71028e-19
cc_118 N_NET21_c_169_n N_Z_c_225_n 7.69306e-19
*
.ends
*
*
.subckt OR2_HPNW12 A B Y VDD VSS
xgate (VSS VDD B A Y) G3_OR2_N3
.ends
*
* File: G4_XNOR2_N3.pex.netlist
* Created: Sun Apr 10 19:31:19 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XNOR2_N3_VDD 2 5 9 12 14 16 32 42 43 45 54 59 66 68 69 70 73 75 76
+ 79 81 85 89 91 93 98 99 100 103 109 114 123 Vss
c102 123 Vss 0.00998345f
c103 114 Vss 0.00466671f
c104 109 Vss 0.00477251f
c105 101 Vss 8.67375e-19
c106 100 Vss 2.39889e-19
c107 99 Vss 4.52364e-19
c108 98 Vss 0.00591503f
c109 93 Vss 0.00301333f
c110 91 Vss 0.0106867f
c111 89 Vss 0.0015063f
c112 85 Vss 6.60056e-19
c113 81 Vss 0.0046084f
c114 79 Vss 0.00109211f
c115 76 Vss 8.68689e-19
c116 75 Vss 0.00224943f
c117 73 Vss 0.00191294f
c118 70 Vss 8.64616e-19
c119 69 Vss 0.00566667f
c120 68 Vss 0.0107726f
c121 66 Vss 0.00280898f
c122 59 Vss 0.00679236f
c123 54 Vss 0.010135f
c124 45 Vss 1.08186e-19
c125 43 Vss 0.0351405f
c126 42 Vss 0.100973f
c127 33 Vss 0.0359366f
c128 32 Vss 0.100971f
c129 14 Vss 0.00143493f
c130 9 Vss 0.377348f
c131 5 Vss 0.379154f
r132 98 103 0.326018
r133 97 98 5.54325
r134 95 123 1.16709
r135 93 97 0.655813
r136 93 95 1.82344
r137 92 101 0.494161
r138 91 103 0.326018
r139 91 92 13.0037
r140 87 101 0.128424
r141 87 89 6.16843
r142 85 114 1.16709
r143 83 85 2.16729
r144 82 100 0.494161
r145 81 101 0.494161
r146 81 82 7.46046
r147 79 109 1.16709
r148 77 100 0.128424
r149 77 79 2.16729
r150 75 100 0.494161
r151 75 76 4.37625
r152 71 99 0.0828784
r153 71 73 1.82344
r154 69 83 0.652036
r155 69 70 10.1279
r156 68 76 0.652036
r157 67 99 0.551426
r158 67 68 17.4633
r159 66 99 0.551426
r160 65 70 0.652036
r161 65 66 5.50157
r162 63 123 0.05
r163 59 89 1.16709
r164 54 73 1.16709
r165 45 114 0.0476429
r166 43 45 1.45875
r167 42 46 0.652036
r168 42 45 1.45875
r169 39 43 0.652036
r170 35 109 0.0476429
r171 33 35 1.45875
r172 32 36 0.652036
r173 32 35 1.45875
r174 29 33 0.652036
r175 16 63 0.123773
r176 14 59 0.123773
r177 12 59 0.123773
r178 9 46 5.1348
r179 9 39 5.1348
r180 5 36 5.1348
r181 5 29 5.1348
r182 2 54 0.123773
.ends

.subckt PM_G4_XNOR2_N3_VSS 3 6 8 11 14 16 32 33 42 43 54 59 63 66 71 76 81 87 96
+ 101 114 116 117 118 123 124 129 137 142 143 144 146 Vss
c85 144 Vss 3.75522e-19
c86 143 Vss 4.28045e-19
c87 142 Vss 0.0047306f
c88 137 Vss 0.00122865f
c89 129 Vss 0.0130341f
c90 124 Vss 8.2479e-19
c91 123 Vss 0.00464476f
c92 118 Vss 8.46757e-19
c93 117 Vss 0.00174235f
c94 116 Vss 0.00202335f
c95 114 Vss 0.00643502f
c96 101 Vss 0.00391102f
c97 96 Vss 0.00421609f
c98 87 Vss 2.60675e-19
c99 81 Vss 0.00257188f
c100 76 Vss 7.28175e-19
c101 71 Vss 0.00117992f
c102 66 Vss 0.00174295f
c103 63 Vss 0.00812841f
c104 59 Vss 0.00683037f
c105 54 Vss 0.00816767f
c106 43 Vss 0.0342891f
c107 42 Vss 0.100071f
c108 33 Vss 0.0350852f
c109 32 Vss 0.0990713f
c110 14 Vss 0.00143493f
c111 11 Vss 0.378924f
c112 3 Vss 0.378636f
r113 142 146 0.349767
r114 141 142 5.50157
r115 137 146 0.306046
r116 130 144 0.494161
r117 129 141 0.652036
r118 125 144 0.128424
r119 123 133 0.652036
r120 123 124 10.1279
r121 119 143 0.0828784
r122 117 144 0.494161
r123 117 118 4.37625
r124 116 124 0.652036
r125 115 143 0.551426
r126 115 116 5.50157
r127 114 143 0.551426
r128 113 118 0.652036
r129 113 114 17.4633
r130 87 137 1.82344
r131 81 129 13.5872
r132 81 130 8.04396
r133 81 84 6.71025
r134 76 101 1.16709
r135 76 133 2.16729
r136 71 96 1.16709
r137 71 125 2.16729
r138 66 119 1.82344
r139 63 87 1.16709
r140 59 84 1.16709
r141 54 66 1.16709
r142 45 101 0.0476429
r143 43 45 1.45875
r144 42 46 0.652036
r145 42 45 1.45875
r146 39 43 0.652036
r147 35 96 0.0476429
r148 33 35 1.45875
r149 32 36 0.652036
r150 32 35 1.45875
r151 29 33 0.652036
r152 16 63 0.123773
r153 14 59 0.123773
r154 11 46 5.1348
r155 11 39 5.1348
r156 8 59 0.123773
r157 6 54 0.123773
r158 3 36 5.1348
r159 3 29 5.1348
.ends

.subckt PM_G4_XNOR2_N3_A 2 4 7 10 21 24 28 39 48 54 57 62 67 72 77 85 Vss
c54 85 Vss 5.19577e-19
c55 77 Vss 0.00107525f
c56 72 Vss 0.00526551f
c57 67 Vss 0.00394354f
c58 62 Vss 0.00276499f
c59 57 Vss 0.00595775f
c60 54 Vss 8.99321e-19
c61 48 Vss 0.126065f
c62 43 Vss 0.0296855f
c63 39 Vss 4.49964e-19
c64 28 Vss 0.152703f
c65 24 Vss 8.95828e-20
c66 21 Vss 0.173355f
c67 18 Vss 0.180502f
c68 16 Vss 0.0247918f
c69 10 Vss 0.176514f
c70 7 Vss 0.433917f
c71 4 Vss 0.193054f
r72 81 85 0.653045
r73 62 77 1.16709
r74 62 85 4.9014
r75 57 72 1.16709
r76 57 81 11.3366
r77 51 67 1.16709
r78 51 54 0.0364688
r79 47 72 0.0238214
r80 47 48 2.334
r81 44 47 2.20433
r82 39 77 0.404964
r83 33 48 0.00605528
r84 31 44 0.00605528
r85 29 43 0.494161
r86 28 30 0.652036
r87 28 29 4.84305
r88 25 43 0.128424
r89 24 67 0.0476429
r90 22 24 0.326018
r91 22 24 0.1167
r92 21 43 0.494161
r93 21 24 6.7686
r94 18 67 0.357321
r95 16 24 0.326018
r96 16 18 0.40845
r97 10 39 4.60965
r98 7 33 5.1348
r99 7 31 5.1348
r100 7 30 5.1348
r101 4 25 5.1348
r102 2 18 4.72635
.ends

.subckt PM_G4_XNOR2_N3_NET1 2 4 7 10 30 31 35 41 44 49 58 66 Vss
c34 66 Vss 2.27666e-19
c35 58 Vss 0.0070279f
c36 49 Vss 0.00633509f
c37 44 Vss 0.0011111f
c38 41 Vss 0.00508953f
c39 35 Vss 0.103132f
c40 31 Vss 0.128995f
c41 30 Vss 9.4155e-20
c42 10 Vss 0.290846f
c43 7 Vss 0.485246f
c44 4 Vss 0.00143493f
r45 62 66 0.653045
r46 49 58 1.16709
r47 49 66 12.9148
r48 44 62 3.37596
r49 41 44 1.16709
r50 33 35 1.70187
r51 30 58 0.0238214
r52 30 31 2.20433
r53 27 30 2.334
r54 25 35 0.17282
r55 24 31 0.00605528
r56 21 33 0.17282
r57 18 27 0.00605528
r58 10 21 8.34405
r59 7 25 7.002
r60 7 24 5.1348
r61 7 18 5.1348
r62 4 41 0.123773
r63 2 41 0.123773
.ends

.subckt PM_G4_XNOR2_N3_NET3 2 4 6 9 21 22 33 39 42 47 56 74 Vss
c47 74 Vss 3.98722e-19
c48 56 Vss 0.00391617f
c49 47 Vss 0.00744607f
c50 42 Vss 0.00230693f
c51 39 Vss 0.00508953f
c52 33 Vss 0.12548f
c53 22 Vss 0.0328697f
c54 21 Vss 0.175168f
c55 9 Vss 0.574903f
c56 6 Vss 0.200347f
c57 4 Vss 0.00143493f
r58 70 74 0.660011
r59 47 56 1.16709
r60 47 74 11.3611
r61 42 70 3.29261
r62 39 42 1.16709
r63 32 56 0.0238214
r64 32 33 2.26917
r65 29 32 2.26917
r66 26 33 0.00605528
r67 24 29 0.00605528
r68 21 23 0.652036
r69 21 22 4.84305
r70 18 22 0.652036
r71 9 26 5.1348
r72 9 24 5.1348
r73 9 23 10.0362
r74 6 18 5.54325
r75 4 39 0.123773
r76 2 39 0.123773
.ends

.subckt PM_G4_XNOR2_N3_B 2 4 7 10 19 20 28 31 33 37 38 48 52 55 58 61 Vss
c34 61 Vss 0.0283565f
c35 55 Vss 0.00145453f
c36 52 Vss 0.136463f
c37 48 Vss 0.0595773f
c38 38 Vss 0.0333783f
c39 37 Vss 0.0913542f
c40 33 Vss 0.0446983f
c41 31 Vss 8.50018e-20
c42 28 Vss 0.0899906f
c43 20 Vss 0.0348606f
c44 19 Vss 0.173355f
c45 10 Vss 0.264298f
c46 7 Vss 0.429172f
c47 4 Vss 0.180506f
c48 2 Vss 0.192541f
r49 55 61 1.16709
r50 55 58 0.0416786
r51 50 52 4.53833
r52 47 48 1.167
r53 42 52 0.00605528
r54 37 39 0.652036
r55 37 38 2.04225
r56 35 48 0.0685365
r57 34 50 0.00605528
r58 33 38 0.652036
r59 32 47 0.0685365
r60 32 33 1.69215
r61 31 61 0.181909
r62 29 61 0.494161
r63 29 31 0.1167
r64 28 47 0.5835
r65 28 31 3.55935
r66 23 61 0.128424
r67 23 61 0.40845
r68 22 61 0.181909
r69 20 22 6.7686
r70 19 61 0.494161
r71 19 22 0.1167
r72 16 20 0.652036
r73 10 39 7.5855
r74 7 42 5.1348
r75 7 35 5.1348
r76 7 34 5.1348
r77 4 61 4.72635
r78 2 16 5.1348
.ends

.subckt PM_G4_XNOR2_N3_Z 2 4 6 8 23 27 30 33 Vss
c28 30 Vss 0.0035978f
c29 27 Vss 0.00609752f
c30 23 Vss 0.00569635f
c31 8 Vss 0.00143493f
c32 6 Vss 0.00143493f
r33 33 35 5.29318
r34 30 33 6.66857
r35 27 35 1.16709
r36 23 30 1.16709
r37 8 27 0.123773
r38 6 23 0.123773
r39 4 27 0.123773
r40 2 23 0.123773
.ends

.subckt G4_XNOR2_N3  VDD VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* VDD	VDD
XI20.X0 N_NET1_XI20.X0_D N_VSS_XI20.X0_PGD N_B_XI20.X0_CG N_VSS_XI20.X0_PGD
+ N_VDD_XI20.X0_S TIGFET_HPNW12
XI24.X0 N_NET3_XI24.X0_D N_VDD_XI24.X0_PGD N_A_XI24.X0_CG N_VDD_XI24.X0_PGD
+ N_VSS_XI24.X0_S TIGFET_HPNW12
XI22.X0 N_NET1_XI22.X0_D N_VDD_XI22.X0_PGD N_B_XI22.X0_CG N_VDD_XI22.X0_PGD
+ N_VSS_XI22.X0_S TIGFET_HPNW12
XI26.X0 N_NET3_XI26.X0_D N_VSS_XI26.X0_PGD N_A_XI26.X0_CG N_VSS_XI26.X0_PGD
+ N_VDD_XI26.X0_S TIGFET_HPNW12
XI21.X0 N_Z_XI21.X0_D N_B_XI21.X0_PGD N_NET3_XI21.X0_CG N_B_XI21.X0_PGD
+ N_VSS_XI21.X0_S TIGFET_HPNW12
XI25.X0 N_Z_XI25.X0_D N_A_XI25.X0_PGD N_B_XI25.X0_CG N_A_XI25.X0_PGD
+ N_VDD_XI25.X0_S TIGFET_HPNW12
XI23.X0 N_Z_XI23.X0_D N_NET1_XI23.X0_PGD N_A_XI23.X0_CG N_NET1_XI23.X0_PGD
+ N_VSS_XI23.X0_S TIGFET_HPNW12
XI27.X0 N_Z_XI27.X0_D N_NET3_XI27.X0_PGD N_NET1_XI27.X0_CG N_NET3_XI27.X0_PGD
+ N_VDD_XI27.X0_S TIGFET_HPNW12
*
x_PM_G4_XNOR2_N3_VDD N_VDD_XI20.X0_S N_VDD_XI24.X0_PGD N_VDD_XI22.X0_PGD
+ N_VDD_XI26.X0_S N_VDD_XI25.X0_S N_VDD_XI27.X0_S N_VDD_c_9_p N_VDD_c_23_p
+ N_VDD_c_5_p N_VDD_c_89_p N_VDD_c_64_p N_VDD_c_11_p N_VDD_c_7_p N_VDD_c_12_p
+ N_VDD_c_6_p N_VDD_c_39_p N_VDD_c_13_p N_VDD_c_14_p N_VDD_c_43_p N_VDD_c_19_p
+ N_VDD_c_10_p N_VDD_c_17_p N_VDD_c_4_p N_VDD_c_53_p N_VDD_c_45_p N_VDD_c_59_p
+ N_VDD_c_36_p N_VDD_c_42_p VDD N_VDD_c_22_p N_VDD_c_18_p N_VDD_c_97_p Vss
+ PM_G4_XNOR2_N3_VDD
x_PM_G4_XNOR2_N3_VSS N_VSS_XI20.X0_PGD N_VSS_XI24.X0_S N_VSS_XI22.X0_S
+ N_VSS_XI26.X0_PGD N_VSS_XI21.X0_S N_VSS_XI23.X0_S N_VSS_c_107_n N_VSS_c_109_n
+ N_VSS_c_154_p N_VSS_c_111_n N_VSS_c_170_p N_VSS_c_113_n N_VSS_c_181_p
+ N_VSS_c_114_n N_VSS_c_117_n N_VSS_c_121_n N_VSS_c_125_n N_VSS_c_183_p
+ N_VSS_c_129_n N_VSS_c_133_n N_VSS_c_136_n N_VSS_c_139_n N_VSS_c_140_n
+ N_VSS_c_141_n N_VSS_c_142_n N_VSS_c_145_n N_VSS_c_146_n N_VSS_c_147_n
+ N_VSS_c_165_p N_VSS_c_148_n N_VSS_c_149_n VSS Vss PM_G4_XNOR2_N3_VSS
x_PM_G4_XNOR2_N3_A N_A_XI24.X0_CG N_A_XI26.X0_CG N_A_XI25.X0_PGD N_A_XI23.X0_CG
+ N_A_c_189_n N_A_c_191_n N_A_c_192_n N_A_c_215_p N_A_c_193_n A N_A_c_197_n
+ N_A_c_216_p N_A_c_200_n N_A_c_202_n N_A_c_214_p N_A_c_212_n Vss
+ PM_G4_XNOR2_N3_A
x_PM_G4_XNOR2_N3_NET1 N_NET1_XI20.X0_D N_NET1_XI22.X0_D N_NET1_XI23.X0_PGD
+ N_NET1_XI27.X0_CG N_NET1_c_263_n N_NET1_c_274_p N_NET1_c_267_p N_NET1_c_242_n
+ N_NET1_c_245_n N_NET1_c_249_n N_NET1_c_257_n N_NET1_c_258_n Vss
+ PM_G4_XNOR2_N3_NET1
x_PM_G4_XNOR2_N3_NET3 N_NET3_XI24.X0_D N_NET3_XI26.X0_D N_NET3_XI21.X0_CG
+ N_NET3_XI27.X0_PGD N_NET3_c_298_n N_NET3_c_314_p N_NET3_c_277_n N_NET3_c_278_n
+ N_NET3_c_279_n N_NET3_c_282_n N_NET3_c_285_n N_NET3_c_287_n Vss
+ PM_G4_XNOR2_N3_NET3
x_PM_G4_XNOR2_N3_B N_B_XI20.X0_CG N_B_XI22.X0_CG N_B_XI21.X0_PGD N_B_XI25.X0_CG
+ N_B_c_325_n N_B_c_338_n N_B_c_327_n N_B_c_328_n N_B_c_351_n N_B_c_347_n
+ N_B_c_340_n N_B_c_341_n N_B_c_329_n N_B_c_330_n B N_B_c_331_n Vss
+ PM_G4_XNOR2_N3_B
x_PM_G4_XNOR2_N3_Z N_Z_XI21.X0_D N_Z_XI25.X0_D N_Z_XI23.X0_D N_Z_XI27.X0_D
+ N_Z_c_367_n N_Z_c_357_n N_Z_c_362_n Z Vss PM_G4_XNOR2_N3_Z
cc_1 N_VDD_XI24.X0_PGD N_VSS_XI20.X0_PGD 2.9783e-19
cc_2 N_VDD_XI22.X0_PGD N_VSS_XI20.X0_PGD 0.0019598f
cc_3 N_VDD_XI24.X0_PGD N_VSS_XI26.X0_PGD 0.0019593f
cc_4 N_VDD_c_4_p N_VSS_XI26.X0_PGD 2.21956e-19
cc_5 N_VDD_c_5_p N_VSS_c_107_n 0.0019598f
cc_6 N_VDD_c_6_p N_VSS_c_107_n 3.89167e-19
cc_7 N_VDD_c_7_p N_VSS_c_109_n 3.80615e-19
cc_8 N_VDD_c_6_p N_VSS_c_109_n 3.89167e-19
cc_9 N_VDD_c_9_p N_VSS_c_111_n 0.0019593f
cc_10 N_VDD_c_10_p N_VSS_c_111_n 3.89167e-19
cc_11 N_VDD_c_11_p N_VSS_c_113_n 3.47417e-19
cc_12 N_VDD_c_12_p N_VSS_c_114_n 0.00187494f
cc_13 N_VDD_c_13_p N_VSS_c_114_n 4.32036e-19
cc_14 N_VDD_c_14_p N_VSS_c_114_n 3.5277e-19
cc_15 N_VDD_c_7_p N_VSS_c_117_n 4.35319e-19
cc_16 N_VDD_c_6_p N_VSS_c_117_n 0.00161703f
cc_17 N_VDD_c_17_p N_VSS_c_117_n 8.66259e-19
cc_18 N_VDD_c_18_p N_VSS_c_117_n 3.48267e-19
cc_19 N_VDD_c_19_p N_VSS_c_121_n 9.53113e-19
cc_20 N_VDD_c_10_p N_VSS_c_121_n 0.00161703f
cc_21 N_VDD_c_4_p N_VSS_c_121_n 0.00227183f
cc_22 N_VDD_c_22_p N_VSS_c_121_n 3.48267e-19
cc_23 N_VDD_c_23_p N_VSS_c_125_n 2.36481e-19
cc_24 N_VDD_c_6_p N_VSS_c_125_n 0.00538298f
cc_25 N_VDD_c_4_p N_VSS_c_125_n 2.5578e-19
cc_26 N_VDD_c_18_p N_VSS_c_125_n 9.58524e-19
cc_27 N_VDD_c_7_p N_VSS_c_129_n 3.66936e-19
cc_28 N_VDD_c_6_p N_VSS_c_129_n 2.26455e-19
cc_29 N_VDD_c_17_p N_VSS_c_129_n 3.99794e-19
cc_30 N_VDD_c_18_p N_VSS_c_129_n 6.489e-19
cc_31 N_VDD_c_10_p N_VSS_c_133_n 2.26455e-19
cc_32 N_VDD_c_4_p N_VSS_c_133_n 9.55322e-19
cc_33 N_VDD_c_22_p N_VSS_c_133_n 6.46219e-19
cc_34 N_VDD_c_7_p N_VSS_c_136_n 0.00378845f
cc_35 N_VDD_c_12_p N_VSS_c_136_n 0.00917884f
cc_36 N_VDD_c_36_p N_VSS_c_136_n 0.0010706f
cc_37 N_VDD_c_12_p N_VSS_c_139_n 0.00404533f
cc_38 N_VDD_c_6_p N_VSS_c_140_n 0.00348469f
cc_39 N_VDD_c_39_p N_VSS_c_141_n 0.00107963f
cc_40 N_VDD_c_14_p N_VSS_c_142_n 0.00356332f
cc_41 N_VDD_c_10_p N_VSS_c_142_n 0.00615517f
cc_42 N_VDD_c_42_p N_VSS_c_142_n 9.37919e-19
cc_43 N_VDD_c_43_p N_VSS_c_145_n 0.00106367f
cc_44 N_VDD_c_6_p N_VSS_c_146_n 0.00468936f
cc_45 N_VDD_c_45_p N_VSS_c_147_n 9.00324e-19
cc_46 N_VDD_c_12_p N_VSS_c_148_n 9.16632e-19
cc_47 N_VDD_c_6_p N_VSS_c_149_n 7.74609e-19
cc_48 N_VDD_c_4_p N_A_XI25.X0_PGD 2.05446e-19
cc_49 N_VDD_XI24.X0_PGD N_A_c_189_n 4.09718e-19
cc_50 N_VDD_XI22.X0_PGD N_A_c_189_n 2.22577e-19
cc_51 N_VDD_c_22_p N_A_c_191_n 5.33384e-19
cc_52 N_VDD_XI22.X0_PGD N_A_c_192_n 2.22577e-19
cc_53 N_VDD_c_53_p N_A_c_193_n 6.08999e-19
cc_54 N_VDD_c_12_p A 5.04211e-19
cc_55 N_VDD_c_19_p A 2.95248e-19
cc_56 N_VDD_c_22_p A 2.15082e-19
cc_57 N_VDD_c_4_p N_A_c_197_n 0.00289813f
cc_58 N_VDD_c_53_p N_A_c_197_n 0.00191817f
cc_59 N_VDD_c_59_p N_A_c_197_n 3.22661e-19
cc_60 N_VDD_c_12_p N_A_c_200_n 6.25289e-19
cc_61 N_VDD_c_19_p N_A_c_200_n 2.28697e-19
cc_62 N_VDD_c_4_p N_A_c_202_n 9.84209e-19
cc_63 N_VDD_c_53_p N_A_c_202_n 2.68554e-19
cc_64 N_VDD_c_64_p N_NET1_c_242_n 3.43419e-19
cc_65 N_VDD_c_6_p N_NET1_c_242_n 2.74986e-19
cc_66 N_VDD_c_13_p N_NET1_c_242_n 3.72199e-19
cc_67 N_VDD_c_64_p N_NET1_c_245_n 3.48267e-19
cc_68 N_VDD_c_7_p N_NET1_c_245_n 2.34601e-19
cc_69 N_VDD_c_6_p N_NET1_c_245_n 2.9533e-19
cc_70 N_VDD_c_13_p N_NET1_c_245_n 5.226e-19
cc_71 N_VDD_c_17_p N_NET1_c_249_n 0.00122163f
cc_72 N_VDD_c_59_p N_NET3_XI27.X0_PGD 4.14305e-19
cc_73 N_VDD_c_53_p N_NET3_c_277_n 8.42825e-19
cc_74 N_VDD_c_11_p N_NET3_c_278_n 3.43419e-19
cc_75 N_VDD_c_11_p N_NET3_c_279_n 3.48267e-19
cc_76 N_VDD_c_10_p N_NET3_c_279_n 3.21336e-19
cc_77 N_VDD_c_4_p N_NET3_c_279_n 0.00123864f
cc_78 N_VDD_c_4_p N_NET3_c_282_n 0.00123016f
cc_79 N_VDD_c_53_p N_NET3_c_282_n 0.00291325f
cc_80 N_VDD_c_59_p N_NET3_c_282_n 7.77543e-19
cc_81 N_VDD_c_53_p N_NET3_c_285_n 0.00118178f
cc_82 N_VDD_c_59_p N_NET3_c_285_n 3.66936e-19
cc_83 N_VDD_c_19_p N_NET3_c_287_n 3.02266e-19
cc_84 N_VDD_c_12_p N_B_XI20.X0_CG 3.50093e-19
cc_85 N_VDD_XI22.X0_PGD N_B_XI21.X0_PGD 0.00190378f
cc_86 N_VDD_XI24.X0_PGD N_B_c_325_n 2.22577e-19
cc_87 N_VDD_XI22.X0_PGD N_B_c_325_n 4.09718e-19
cc_88 N_VDD_XI22.X0_PGD N_B_c_327_n 4.09718e-19
cc_89 N_VDD_c_89_p N_B_c_328_n 5.7019e-19
cc_90 N_VDD_c_23_p N_B_c_329_n 0.00168656f
cc_91 N_VDD_c_18_p N_B_c_330_n 2.15082e-19
cc_92 N_VDD_c_17_p N_B_c_331_n 2.26584e-19
cc_93 N_VDD_c_11_p N_Z_c_357_n 3.43419e-19
cc_94 N_VDD_c_4_p N_Z_c_357_n 3.48267e-19
cc_95 N_VDD_c_53_p N_Z_c_357_n 2.74986e-19
cc_96 N_VDD_c_45_p N_Z_c_357_n 3.72199e-19
cc_97 N_VDD_c_97_p N_Z_c_357_n 3.43419e-19
cc_98 N_VDD_c_11_p N_Z_c_362_n 3.48267e-19
cc_99 N_VDD_c_4_p N_Z_c_362_n 4.85404e-19
cc_100 N_VDD_c_53_p N_Z_c_362_n 4.9751e-19
cc_101 N_VDD_c_45_p N_Z_c_362_n 8.21216e-19
cc_102 N_VDD_c_97_p N_Z_c_362_n 3.48267e-19
cc_103 N_VSS_XI26.X0_PGD N_A_XI25.X0_PGD 0.00164979f
cc_104 N_VSS_XI20.X0_PGD N_A_c_189_n 2.22577e-19
cc_105 N_VSS_XI26.X0_PGD N_A_c_189_n 4.09718e-19
cc_106 N_VSS_XI26.X0_PGD N_A_c_192_n 4.09718e-19
cc_107 N_VSS_c_154_p N_A_c_193_n 0.00164979f
cc_108 N_VSS_c_121_n N_A_c_197_n 3.87149e-19
cc_109 N_VSS_c_136_n N_A_c_197_n 6.21456e-19
cc_110 N_VSS_c_133_n N_A_c_202_n 6.52904e-19
cc_111 N_VSS_c_146_n N_A_c_212_n 5.04853e-19
cc_112 N_VSS_c_113_n N_NET1_c_242_n 3.43419e-19
cc_113 N_VSS_c_125_n N_NET1_c_242_n 3.48267e-19
cc_114 N_VSS_c_113_n N_NET1_c_245_n 3.48267e-19
cc_115 N_VSS_c_125_n N_NET1_c_245_n 0.00164479f
cc_116 N_VSS_c_125_n N_NET1_c_249_n 0.00162978f
cc_117 N_VSS_c_146_n N_NET1_c_249_n 0.0181004f
cc_118 N_VSS_c_165_p N_NET1_c_249_n 0.00121213f
cc_119 N_VSS_c_125_n N_NET1_c_257_n 2.78343e-19
cc_120 N_VSS_c_117_n N_NET1_c_258_n 0.00198862f
cc_121 N_VSS_c_136_n N_NET1_c_258_n 0.00136675f
cc_122 N_VSS_c_146_n N_NET1_c_258_n 0.00168829f
cc_123 N_VSS_c_170_p N_NET3_c_278_n 3.43419e-19
cc_124 N_VSS_c_170_p N_NET3_c_279_n 3.48267e-19
cc_125 N_VSS_c_114_n N_NET3_c_279_n 0.0011211f
cc_126 N_VSS_c_139_n N_NET3_c_279_n 6.33709e-19
cc_127 N_VSS_c_121_n N_NET3_c_282_n 0.00131985f
cc_128 N_VSS_c_142_n N_NET3_c_287_n 4.84133e-19
cc_129 N_VSS_XI20.X0_PGD N_B_c_325_n 4.09718e-19
cc_130 N_VSS_XI26.X0_PGD N_B_c_325_n 2.22577e-19
cc_131 N_VSS_XI26.X0_PGD N_B_c_327_n 2.22577e-19
cc_132 N_VSS_c_125_n N_B_c_329_n 2.44335e-19
cc_133 N_VSS_c_113_n N_Z_c_367_n 3.43419e-19
cc_134 N_VSS_c_181_p N_Z_c_367_n 3.43419e-19
cc_135 N_VSS_c_125_n N_Z_c_367_n 3.48267e-19
cc_136 N_VSS_c_183_p N_Z_c_367_n 3.48267e-19
cc_137 N_VSS_c_113_n N_Z_c_362_n 3.48267e-19
cc_138 N_VSS_c_181_p N_Z_c_362_n 3.48267e-19
cc_139 N_VSS_c_125_n N_Z_c_362_n 8.69457e-19
cc_140 N_VSS_c_183_p N_Z_c_362_n 5.71987e-19
cc_141 N_A_XI23.X0_CG N_NET1_XI23.X0_PGD 5.00154e-19
cc_142 N_A_c_214_p N_NET1_XI23.X0_PGD 0.0013363f
cc_143 N_A_c_215_p N_NET1_c_263_n 5.8445e-19
cc_144 N_A_c_216_p N_NET1_c_249_n 0.0020999f
cc_145 N_A_c_212_n N_NET1_c_249_n 6.74055e-19
cc_146 N_A_c_214_p N_NET3_XI21.X0_CG 2.18475e-19
cc_147 N_A_XI25.X0_PGD N_NET3_XI27.X0_PGD 0.00173934f
cc_148 N_A_c_192_n N_NET3_XI27.X0_PGD 3.14428e-19
cc_149 N_A_c_214_p N_NET3_XI27.X0_PGD 4.34237e-19
cc_150 N_A_XI25.X0_PGD N_NET3_c_298_n 4.64512e-19
cc_151 N_A_c_193_n N_NET3_c_277_n 0.00173934f
cc_152 N_A_c_189_n N_NET3_c_278_n 6.35441e-19
cc_153 N_A_c_197_n N_NET3_c_279_n 0.00122226f
cc_154 N_A_c_197_n N_NET3_c_282_n 0.00256249f
cc_155 N_A_c_216_p N_NET3_c_282_n 0.00124966f
cc_156 N_A_c_202_n N_NET3_c_282_n 3.44698e-19
cc_157 N_A_c_197_n N_NET3_c_285_n 3.44698e-19
cc_158 N_A_c_202_n N_NET3_c_285_n 6.70706e-19
cc_159 N_A_c_192_n N_B_XI25.X0_CG 0.003858f
cc_160 N_A_c_189_n N_B_c_325_n 0.00503082f
cc_161 N_A_c_200_n N_B_c_338_n 7.5077e-19
cc_162 N_A_c_192_n N_B_c_327_n 0.00270268f
cc_163 N_A_c_192_n N_B_c_340_n 0.00358164f
cc_164 N_A_c_192_n N_B_c_341_n 2.04018e-19
cc_165 N_A_c_212_n N_B_c_330_n 2.24721e-19
cc_166 N_A_c_189_n N_B_c_331_n 8.36919e-19
cc_167 N_A_c_197_n N_Z_c_362_n 0.00453915f
cc_168 N_A_c_216_p N_Z_c_362_n 0.00285282f
cc_169 N_A_c_214_p N_Z_c_362_n 9.79999e-19
cc_170 N_NET1_XI23.X0_PGD N_NET3_XI21.X0_CG 3.25363e-19
cc_171 N_NET1_c_267_p N_NET3_XI27.X0_PGD 0.00866857f
cc_172 N_NET1_XI23.X0_PGD N_NET3_c_298_n 0.00335065f
cc_173 N_NET1_c_242_n N_NET3_c_278_n 2.56771e-19
cc_174 N_NET1_XI23.X0_PGD N_B_XI21.X0_PGD 0.00216073f
cc_175 N_NET1_XI27.X0_CG N_B_XI25.X0_CG 2.72501e-19
cc_176 N_NET1_c_242_n N_B_c_325_n 6.35441e-19
cc_177 N_NET1_c_267_p N_B_c_347_n 2.72501e-19
cc_178 N_NET1_c_274_p N_B_c_329_n 0.00193498f
cc_179 N_NET1_c_249_n N_Z_c_362_n 3.17674e-19
cc_180 N_NET3_XI21.X0_CG N_B_XI21.X0_PGD 0.00200964f
cc_181 N_NET3_c_298_n N_B_XI21.X0_PGD 0.00163867f
cc_182 N_NET3_XI27.X0_PGD N_B_c_351_n 3.23792e-19
cc_183 N_NET3_c_314_p N_B_c_351_n 5.75226e-19
cc_184 N_NET3_XI27.X0_PGD N_B_c_347_n 0.00310335f
cc_185 N_NET3_c_314_p N_B_c_347_n 0.00201276f
cc_186 N_NET3_c_314_p N_B_c_341_n 0.00200964f
cc_187 N_NET3_c_298_n N_Z_c_367_n 6.58359e-19
cc_188 N_NET3_c_298_n N_Z_c_357_n 2.51847e-19
cc_189 N_NET3_XI27.X0_PGD N_Z_c_362_n 0.00129454f
cc_190 N_NET3_c_298_n N_Z_c_362_n 2.39178e-19
cc_191 N_NET3_c_282_n N_Z_c_362_n 2.33494e-19
cc_192 N_B_c_347_n N_Z_c_362_n 9.47639e-19
*
.ends
*
*
.subckt XNOR2_HPNW12 A B Y VDD VSS
xgate (VDD VSS A B Y) G4_XNOR2_N3
.ends
*
* File: G5_XNOR3_N3.pex.netlist
* Created: Mon Mar 28 16:13:50 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XNOR3_N3_VDD 2 5 9 12 14 17 34 35 44 45 54 55 65 69 74 77 79 80 81
+ 84 86 87 90 93 96 98 102 104 108 112 114 116 117 119 125 134 139 Vss
c113 139 Vss 0.0048986f
c114 134 Vss 0.00495479f
c115 125 Vss 0.00563771f
c116 117 Vss 2.39889e-19
c117 116 Vss 4.92173e-19
c118 115 Vss 5.21614e-19
c119 114 Vss 4.52364e-19
c120 112 Vss 0.0017155f
c121 110 Vss 0.00173699f
c122 108 Vss 6.49327e-19
c123 104 Vss 0.00471178f
c124 102 Vss 0.0010418f
c125 98 Vss 0.00587581f
c126 96 Vss 0.00147489f
c127 93 Vss 0.00334883f
c128 90 Vss 0.00547221f
c129 87 Vss 8.67855e-19
c130 86 Vss 0.00654417f
c131 84 Vss 0.00154142f
c132 81 Vss 8.68392e-19
c133 80 Vss 0.00938293f
c134 79 Vss 0.0116507f
c135 77 Vss 0.00304889f
c136 74 Vss 0.00785043f
c137 69 Vss 0.00836757f
c138 65 Vss 0.00811483f
c139 55 Vss 0.0356247f
c140 54 Vss 0.10084f
c141 45 Vss 0.0356281f
c142 44 Vss 0.101312f
c143 35 Vss 0.0346562f
c144 34 Vss 0.0991017f
c145 17 Vss 0.378772f
c146 9 Vss 0.379175f
c147 5 Vss 0.383323f
r148 110 119 0.326018
r149 110 112 6.16843
r150 108 139 1.16709
r151 106 108 2.16729
r152 105 117 0.494161
r153 104 119 0.326018
r154 104 105 7.46046
r155 102 134 1.16709
r156 100 117 0.128424
r157 100 102 2.16729
r158 99 116 0.494161
r159 98 106 0.652036
r160 98 99 10.3363
r161 94 115 0.0828784
r162 94 96 2.00578
r163 93 116 0.128424
r164 92 115 0.551426
r165 92 93 5.50157
r166 90 125 1.16709
r167 88 115 0.551426
r168 88 90 7.66886
r169 86 116 0.494161
r170 86 87 10.1279
r171 82 114 0.0828784
r172 82 84 1.82344
r173 80 117 0.494161
r174 80 81 15.8795
r175 79 87 0.652036
r176 78 114 0.551426
r177 78 79 18.3386
r178 77 114 0.551426
r179 76 81 0.652036
r180 76 77 5.50157
r181 74 112 1.16709
r182 69 96 1.16709
r183 65 84 1.16709
r184 57 139 0.0476429
r185 55 57 1.45875
r186 54 58 0.652036
r187 54 57 1.45875
r188 51 55 0.652036
r189 47 134 0.0476429
r190 45 47 1.45875
r191 44 48 0.652036
r192 44 47 1.45875
r193 41 45 0.652036
r194 37 125 0.238214
r195 35 37 1.45875
r196 34 38 0.652036
r197 34 37 1.45875
r198 31 35 0.652036
r199 17 58 5.1348
r200 17 51 5.1348
r201 14 74 0.123773
r202 12 69 0.123773
r203 9 48 5.1348
r204 9 41 5.1348
r205 5 38 5.1348
r206 5 31 5.1348
r207 2 65 0.123773
.ends

.subckt PM_G5_XNOR3_N3_C 2 4 6 8 17 20 23 32 37 40 44 47 52 57 84 92 98 Vss
c49 98 Vss 3.10785e-19
c50 92 Vss 0.00560641f
c51 84 Vss 0.00950787f
c52 57 Vss 0.004971f
c53 52 Vss 7.31067e-19
c54 47 Vss 0.00104925f
c55 40 Vss 0.00163759f
c56 37 Vss 0.0082356f
c57 32 Vss 0.00958317f
c58 23 Vss 2.04877e-19
c59 20 Vss 0.221837f
c60 17 Vss 0.180502f
c61 15 Vss 0.0247918f
c62 4 Vss 0.188411f
r63 93 98 0.441572
r64 92 94 0.655813
r65 92 93 9.04425
r66 88 98 0.174814
r67 84 98 0.441572
r68 52 94 3.33429
r69 47 88 3.33429
r70 40 57 1.16709
r71 40 84 22.1365
r72 40 44 0.0833571
r73 37 52 1.16709
r74 32 47 1.16709
r75 23 57 0.0476429
r76 21 23 0.326018
r77 21 23 0.1167
r78 20 24 0.652036
r79 20 23 6.7686
r80 17 57 0.357321
r81 15 23 0.326018
r82 15 17 0.40845
r83 8 37 0.123773
r84 6 32 0.123773
r85 4 24 5.1348
r86 2 17 4.72635
.ends

.subckt PM_G5_XNOR3_N3_VSS 3 6 8 11 15 18 34 37 44 45 54 55 57 66 70 73 78 83 88
+ 93 96 99 108 113 122 124 125 126 131 132 137 149 153 154 155 Vss
c122 155 Vss 3.75522e-19
c123 154 Vss 3.91906e-19
c124 153 Vss 4.4306e-19
c125 149 Vss 3.17876e-19
c126 137 Vss 0.00359616f
c127 132 Vss 8.45126e-19
c128 131 Vss 0.00635332f
c129 126 Vss 8.42189e-19
c130 125 Vss 0.0059194f
c131 124 Vss 0.00452138f
c132 122 Vss 0.00375531f
c133 113 Vss 0.00410359f
c134 108 Vss 0.00419612f
c135 99 Vss 0.00605485f
c136 96 Vss 0.00346991f
c137 93 Vss 0.00310291f
c138 88 Vss 2.34373e-19
c139 83 Vss 0.00134516f
c140 78 Vss 0.0023966f
c141 73 Vss 0.00367309f
c142 70 Vss 0.0100681f
c143 66 Vss 0.00715185f
c144 57 Vss 9.33833e-20
c145 55 Vss 0.0347733f
c146 54 Vss 0.0999406f
c147 45 Vss 0.035088f
c148 44 Vss 0.0994129f
c149 37 Vss 5.39995e-20
c150 35 Vss 0.0349058f
c151 34 Vss 0.100344f
c152 15 Vss 0.379275f
c153 11 Vss 0.379887f
c154 8 Vss 0.00143493f
c155 3 Vss 0.3841f
r156 147 149 0.416786
r157 143 155 0.494161
r158 139 155 0.128424
r159 138 154 0.494161
r160 137 147 0.652036
r161 137 138 7.46046
r162 133 154 0.128424
r163 131 155 0.494161
r164 131 132 15.8795
r165 127 153 0.0828784
r166 125 154 0.494161
r167 125 126 13.0037
r168 124 132 0.652036
r169 123 153 0.551426
r170 123 124 13.8373
r171 122 153 0.551426
r172 121 126 0.652036
r173 121 122 10.0029
r174 96 143 8.04396
r175 93 96 6.75193
r176 88 113 1.16709
r177 88 149 1.7505
r178 83 108 1.16709
r179 83 139 2.16729
r180 78 133 6.16843
r181 73 99 1.16709
r182 73 127 4.33978
r183 70 93 1.16709
r184 66 78 1.16709
r185 57 113 0.0476429
r186 55 57 1.45875
r187 54 58 0.652036
r188 54 57 1.45875
r189 51 55 0.652036
r190 47 108 0.0476429
r191 45 47 1.45875
r192 44 48 0.652036
r193 44 47 1.45875
r194 41 45 0.652036
r195 37 99 0.238214
r196 35 37 1.45875
r197 34 38 0.652036
r198 34 37 1.45875
r199 31 35 0.652036
r200 18 70 0.123773
r201 15 58 5.1348
r202 15 51 5.1348
r203 11 48 5.1348
r204 11 41 5.1348
r205 8 66 0.123773
r206 6 66 0.123773
r207 3 38 5.1348
r208 3 31 5.1348
.ends

.subckt PM_G5_XNOR3_N3_CI 2 4 6 8 23 26 31 34 39 44 79 80 85 91 Vss
c47 91 Vss 2.55674e-19
c48 85 Vss 0.00650738f
c49 80 Vss 3.61784e-19
c50 79 Vss 0.00547357f
c51 44 Vss 7.31067e-19
c52 39 Vss 7.72278e-19
c53 34 Vss 0.00616608f
c54 31 Vss 0.00967911f
c55 26 Vss 0.00811165f
c56 23 Vss 0.00522928f
c57 4 Vss 0.00143493f
r58 86 91 0.441572
r59 85 87 0.655813
r60 85 86 9.04425
r61 81 91 0.174814
r62 79 91 0.441572
r63 79 80 19.1096
r64 75 80 0.655813
r65 44 87 3.33429
r66 39 81 3.33429
r67 34 75 16.1713
r68 31 44 1.16709
r69 26 39 1.16709
r70 23 34 1.16709
r71 8 31 0.123773
r72 6 26 0.123773
r73 4 23 0.123773
r74 2 23 0.123773
.ends

.subckt PM_G5_XNOR3_N3_A 2 4 7 11 24 44 45 49 51 54 56 57 60 65 66 69 74 Vss
c69 74 Vss 0.00565895f
c70 69 Vss 0.00509443f
c71 66 Vss 0.00618081f
c72 65 Vss 7.10913e-19
c73 57 Vss 8.70991e-19
c74 56 Vss 6.16621e-19
c75 54 Vss 0.00573533f
c76 51 Vss 0.00643922f
c77 49 Vss 0.135088f
c78 45 Vss 0.127808f
c79 44 Vss 1.14131e-19
c80 24 Vss 0.217341f
c81 21 Vss 0.18375f
c82 19 Vss 0.0247918f
c83 7 Vss 1.43795f
c84 4 Vss 0.194116f
r85 65 74 1.16709
r86 65 66 0.531835
r87 62 69 1.16709
r88 60 62 0.125036
r89 57 60 0.708536
r90 56 66 10.4613
r91 53 56 0.652036
r92 53 54 10.503
r93 52 57 0.0685365
r94 51 54 0.652036
r95 51 52 10.2113
r96 47 49 4.53833
r97 44 74 0.0238214
r98 44 45 2.26917
r99 41 44 2.26917
r100 36 49 0.00605528
r101 35 45 0.00605528
r102 32 47 0.00605528
r103 31 41 0.00605528
r104 27 69 0.0952857
r105 25 27 0.326018
r106 25 27 0.1167
r107 24 28 0.652036
r108 24 27 6.7686
r109 21 27 0.3335
r110 19 27 0.326018
r111 19 21 0.2334
r112 11 36 5.1348
r113 11 32 5.1348
r114 7 11 17.9718
r115 7 35 5.1348
r116 7 11 17.9718
r117 7 31 5.1348
r118 4 28 5.1348
r119 2 21 4.9014
.ends

.subckt PM_G5_XNOR3_N3_BI 2 4 6 8 16 23 29 32 37 42 51 56 64 65 68 77 82 83 Vss
c67 83 Vss 7.14146e-20
c68 82 Vss 6.9543e-19
c69 77 Vss 9.4202e-19
c70 68 Vss 6.59929e-19
c71 65 Vss 3.58032e-19
c72 64 Vss 0.00251452f
c73 56 Vss 0.00269072f
c74 51 Vss 0.0023082f
c75 42 Vss 0.00171238f
c76 37 Vss 4.65964e-19
c77 32 Vss 0.00208283f
c78 29 Vss 0.00520899f
c79 23 Vss 9.01088e-20
c80 16 Vss 0.166484f
c81 8 Vss 0.166484f
c82 4 Vss 0.00143493f
r83 81 83 0.65409
r84 81 82 3.42052
r85 77 82 0.652979
r86 68 77 2.03284
r87 66 68 2.00057
r88 64 66 0.652036
r89 64 65 13.2121
r90 60 65 0.652036
r91 42 56 1.16709
r92 42 83 2.00578
r93 37 51 1.16709
r94 37 68 0.0416786
r95 32 60 5.62661
r96 29 32 1.16709
r97 23 56 0.50025
r98 16 51 0.50025
r99 8 23 4.37625
r100 6 16 4.37625
r101 4 29 0.123773
r102 2 29 0.123773
.ends

.subckt PM_G5_XNOR3_N3_AI 2 4 7 11 31 37 43 46 51 60 68 Vss
c46 68 Vss 2.68274e-19
c47 60 Vss 0.00659076f
c48 51 Vss 0.00468816f
c49 46 Vss 8.13811e-19
c50 43 Vss 0.00461167f
c51 37 Vss 0.12791f
c52 31 Vss 0.134438f
c53 7 Vss 1.42501f
c54 4 Vss 0.00143493f
r55 64 68 0.655813
r56 51 60 1.16709
r57 51 68 12.0347
r58 46 64 3.33429
r59 43 46 1.16709
r60 36 60 0.0238214
r61 36 37 2.334
r62 33 36 2.20433
r63 29 31 4.53833
r64 26 37 0.00605528
r65 25 31 0.00605528
r66 22 33 0.00605528
r67 21 29 0.00605528
r68 11 26 5.1348
r69 11 22 5.1348
r70 7 11 17.9718
r71 7 25 5.1348
r72 7 11 17.9718
r73 7 21 5.1348
r74 4 43 0.123773
r75 2 43 0.123773
.ends

.subckt PM_G5_XNOR3_N3_B 2 4 6 8 16 17 24 31 41 44 49 54 59 65 69 76 77 Vss
c63 77 Vss 3.11913e-19
c64 76 Vss 9.9238e-19
c65 69 Vss 0.00389578f
c66 65 Vss 0.00255458f
c67 59 Vss 0.00150469f
c68 54 Vss 0.00172736f
c69 49 Vss 0.00131253f
c70 44 Vss 1.53364e-19
c71 41 Vss 3.86756e-19
c72 31 Vss 0.166484f
c73 24 Vss 8.82658e-20
c74 20 Vss 0.0247918f
c75 17 Vss 0.0339179f
c76 16 Vss 0.186033f
c77 6 Vss 0.166669f
c78 4 Vss 0.177261f
c79 2 Vss 0.191454f
r80 76 77 0.655813
r81 75 76 4.04282
r82 69 75 0.653045
r83 59 62 0.35
r84 49 65 1.16709
r85 49 77 2.00578
r86 44 59 1.16709
r87 44 69 2.1395
r88 41 54 1.16709
r89 41 44 10.7364
r90 36 54 0.309679
r91 31 65 0.50025
r92 28 62 0.452607
r93 24 54 0.214393
r94 20 36 0.326018
r95 20 24 0.75855
r96 17 36 6.7686
r97 16 36 0.326018
r98 16 36 0.1167
r99 13 17 0.652036
r100 8 31 4.37625
r101 6 28 4.2012
r102 4 24 4.37625
r103 2 13 5.1348
.ends

.subckt PM_G5_XNOR3_N3_Z 2 4 6 8 23 27 30 33 Vss
c30 30 Vss 0.00380939f
c31 27 Vss 0.00807893f
c32 23 Vss 0.00720799f
c33 8 Vss 0.00143493f
c34 6 Vss 0.00143493f
r35 33 35 6.33514
r36 30 33 6.50186
r37 27 35 1.16709
r38 23 30 1.16709
r39 8 27 0.123773
r40 6 23 0.123773
r41 4 27 0.123773
r42 2 23 0.123773
.ends

.subckt G5_XNOR3_N3  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI22.X0 N_CI_XI22.X0_D N_VSS_XI22.X0_PGD N_C_XI22.X0_CG N_VSS_XI22.X0_PGD
+ N_VDD_XI22.X0_S TIGFET_HPNW12
XI26.X0 N_CI_XI26.X0_D N_VDD_XI26.X0_PGD N_C_XI26.X0_CG N_VDD_XI26.X0_PGD
+ N_VSS_XI26.X0_S TIGFET_HPNW12
XI25.X0 N_BI_XI25.X0_D N_VDD_XI25.X0_PGD N_B_XI25.X0_CG N_VDD_XI25.X0_PGD
+ N_VSS_XI25.X0_S TIGFET_HPNW12
XI21.X0 N_AI_XI21.X0_D N_VSS_XI21.X0_PGD N_A_XI21.X0_CG N_VSS_XI21.X0_PGD
+ N_VDD_XI21.X0_S TIGFET_HPNW12
XI23.X0 N_BI_XI23.X0_D N_VSS_XI23.X0_PGD N_B_XI23.X0_CG N_VSS_XI23.X0_PGD
+ N_VDD_XI23.X0_S TIGFET_HPNW12
XI24.X0 N_AI_XI24.X0_D N_VDD_XI24.X0_PGD N_A_XI24.X0_CG N_VDD_XI24.X0_PGD
+ N_VSS_XI24.X0_S TIGFET_HPNW12
XI31.X0 N_Z_XI31.X0_D N_AI_XI31.X0_PGD N_B_XI31.X0_CG N_AI_XI31.X0_PGD
+ N_C_XI31.X0_S TIGFET_HPNW12
XI27.X0 N_Z_XI27.X0_D N_AI_XI27.X0_PGD N_BI_XI27.X0_CG N_AI_XI27.X0_PGD
+ N_CI_XI27.X0_S TIGFET_HPNW12
XI29.X0 N_Z_XI29.X0_D N_A_XI29.X0_PGD N_BI_XI29.X0_CG N_A_XI29.X0_PGD
+ N_C_XI29.X0_S TIGFET_HPNW12
XI28.X0 N_Z_XI28.X0_D N_A_XI28.X0_PGD N_B_XI28.X0_CG N_A_XI28.X0_PGD
+ N_CI_XI28.X0_S TIGFET_HPNW12
*
x_PM_G5_XNOR3_N3_VDD N_VDD_XI22.X0_S N_VDD_XI26.X0_PGD N_VDD_XI25.X0_PGD
+ N_VDD_XI21.X0_S N_VDD_XI23.X0_S N_VDD_XI24.X0_PGD N_VDD_c_112_p N_VDD_c_19_p
+ N_VDD_c_24_p N_VDD_c_4_p N_VDD_c_102_p N_VDD_c_20_p N_VDD_c_78_p N_VDD_c_103_p
+ N_VDD_c_6_p N_VDD_c_7_p N_VDD_c_13_p N_VDD_c_5_p N_VDD_c_64_p N_VDD_c_29_p
+ N_VDD_c_65_p N_VDD_c_69_p N_VDD_c_30_p N_VDD_c_16_p N_VDD_c_66_p N_VDD_c_21_p
+ N_VDD_c_10_p N_VDD_c_25_p N_VDD_c_37_p N_VDD_c_11_p N_VDD_c_60_p N_VDD_c_68_p
+ N_VDD_c_72_p VDD N_VDD_c_2_p N_VDD_c_42_p N_VDD_c_38_p Vss PM_G5_XNOR3_N3_VDD
x_PM_G5_XNOR3_N3_C N_C_XI22.X0_CG N_C_XI26.X0_CG N_C_XI31.X0_S N_C_XI29.X0_S
+ N_C_c_129_p N_C_c_116_n N_C_c_126_p N_C_c_119_n N_C_c_157_p N_C_c_120_n C
+ N_C_c_127_p N_C_c_159_p N_C_c_122_n N_C_c_123_n N_C_c_143_p N_C_c_148_p Vss
+ PM_G5_XNOR3_N3_C
x_PM_G5_XNOR3_N3_VSS N_VSS_XI22.X0_PGD N_VSS_XI26.X0_S N_VSS_XI25.X0_S
+ N_VSS_XI21.X0_PGD N_VSS_XI23.X0_PGD N_VSS_XI24.X0_S N_VSS_c_170_n
+ N_VSS_c_230_n N_VSS_c_171_n N_VSS_c_173_n N_VSS_c_174_n N_VSS_c_175_n
+ N_VSS_c_281_p N_VSS_c_177_n N_VSS_c_242_p N_VSS_c_178_n N_VSS_c_183_n
+ N_VSS_c_186_n N_VSS_c_190_n N_VSS_c_194_n N_VSS_c_197_n N_VSS_c_198_n
+ N_VSS_c_201_n N_VSS_c_205_n N_VSS_c_209_n N_VSS_c_212_n N_VSS_c_214_n
+ N_VSS_c_215_n N_VSS_c_216_n N_VSS_c_220_n N_VSS_c_221_n VSS N_VSS_c_226_n
+ N_VSS_c_227_n N_VSS_c_228_n Vss PM_G5_XNOR3_N3_VSS
x_PM_G5_XNOR3_N3_CI N_CI_XI22.X0_D N_CI_XI26.X0_D N_CI_XI27.X0_S N_CI_XI28.X0_S
+ N_CI_c_285_n N_CI_c_297_n N_CI_c_326_p N_CI_c_286_n N_CI_c_304_n N_CI_c_328_p
+ N_CI_c_290_n N_CI_c_310_n N_CI_c_313_p N_CI_c_322_p Vss PM_G5_XNOR3_N3_CI
x_PM_G5_XNOR3_N3_A N_A_XI21.X0_CG N_A_XI24.X0_CG N_A_XI29.X0_PGD N_A_XI28.X0_PGD
+ N_A_c_332_n N_A_c_361_p N_A_c_373_p N_A_c_375_p N_A_c_333_n N_A_c_338_n
+ N_A_c_339_n N_A_c_340_n A N_A_c_346_n N_A_c_347_n N_A_c_341_n N_A_c_364_p Vss
+ PM_G5_XNOR3_N3_A
x_PM_G5_XNOR3_N3_BI N_BI_XI25.X0_D N_BI_XI23.X0_D N_BI_XI27.X0_CG
+ N_BI_XI29.X0_CG N_BI_c_432_p N_BI_c_423_n N_BI_c_401_n N_BI_c_403_n
+ N_BI_c_437_p N_BI_c_418_n N_BI_c_433_p N_BI_c_427_n N_BI_c_408_n N_BI_c_416_n
+ N_BI_c_431_n N_BI_c_409_n N_BI_c_458_p N_BI_c_410_n Vss PM_G5_XNOR3_N3_BI
x_PM_G5_XNOR3_N3_AI N_AI_XI21.X0_D N_AI_XI24.X0_D N_AI_XI31.X0_PGD
+ N_AI_XI27.X0_PGD N_AI_c_478_n N_AI_c_469_n N_AI_c_470_n N_AI_c_472_n
+ N_AI_c_476_n N_AI_c_485_n N_AI_c_486_n Vss PM_G5_XNOR3_N3_AI
x_PM_G5_XNOR3_N3_B N_B_XI25.X0_CG N_B_XI23.X0_CG N_B_XI31.X0_CG N_B_XI28.X0_CG
+ N_B_c_515_n N_B_c_516_n N_B_c_522_n N_B_c_532_n B N_B_c_535_n N_B_c_526_n
+ N_B_c_537_n N_B_c_540_n N_B_c_542_n N_B_c_517_n N_B_c_563_n N_B_c_566_n Vss
+ PM_G5_XNOR3_N3_B
x_PM_G5_XNOR3_N3_Z N_Z_XI31.X0_D N_Z_XI27.X0_D N_Z_XI29.X0_D N_Z_XI28.X0_D
+ N_Z_c_577_n N_Z_c_584_n N_Z_c_581_n Z Vss PM_G5_XNOR3_N3_Z
cc_1 N_VDD_XI25.X0_PGD N_C_XI26.X0_CG 0.00111653f
cc_2 N_VDD_c_2_p N_C_XI26.X0_CG 0.00108697f
cc_3 N_VDD_XI26.X0_PGD N_C_c_116_n 4.20258e-19
cc_4 N_VDD_c_4_p N_C_c_116_n 0.00111653f
cc_5 N_VDD_c_5_p N_C_c_116_n 0.00135138f
cc_6 N_VDD_c_6_p N_C_c_119_n 3.43419e-19
cc_7 N_VDD_c_7_p N_C_c_120_n 4.76491e-19
cc_8 N_VDD_c_5_p N_C_c_120_n 0.00161703f
cc_9 N_VDD_c_5_p N_C_c_122_n 2.84771e-19
cc_10 N_VDD_c_10_p N_C_c_123_n 5.71495e-19
cc_11 N_VDD_c_11_p N_C_c_123_n 8.59389e-19
cc_12 N_VDD_XI26.X0_PGD N_VSS_XI22.X0_PGD 0.00200994f
cc_13 N_VDD_c_13_p N_VSS_XI22.X0_PGD 4.18763e-19
cc_14 N_VDD_XI25.X0_PGD N_VSS_XI21.X0_PGD 2.44446e-19
cc_15 N_VDD_XI24.X0_PGD N_VSS_XI21.X0_PGD 0.00200236f
cc_16 N_VDD_c_16_p N_VSS_XI21.X0_PGD 4.15609e-19
cc_17 N_VDD_XI25.X0_PGD N_VSS_XI23.X0_PGD 0.00200584f
cc_18 N_VDD_XI24.X0_PGD N_VSS_XI23.X0_PGD 2.31309e-19
cc_19 N_VDD_c_19_p N_VSS_c_170_n 0.00200994f
cc_20 N_VDD_c_20_p N_VSS_c_171_n 0.00200236f
cc_21 N_VDD_c_21_p N_VSS_c_171_n 3.00203e-19
cc_22 N_VDD_c_21_p N_VSS_c_173_n 3.89167e-19
cc_23 N_VDD_c_11_p N_VSS_c_174_n 2.35465e-19
cc_24 N_VDD_c_24_p N_VSS_c_175_n 0.00200584f
cc_25 N_VDD_c_25_p N_VSS_c_175_n 3.89167e-19
cc_26 N_VDD_c_5_p N_VSS_c_177_n 2.74986e-19
cc_27 N_VDD_c_13_p N_VSS_c_178_n 4.32468e-19
cc_28 N_VDD_c_5_p N_VSS_c_178_n 3.08724e-19
cc_29 N_VDD_c_29_p N_VSS_c_178_n 0.00111881f
cc_30 N_VDD_c_30_p N_VSS_c_178_n 3.98949e-19
cc_31 N_VDD_c_2_p N_VSS_c_178_n 3.48267e-19
cc_32 N_VDD_c_5_p N_VSS_c_183_n 2.9533e-19
cc_33 N_VDD_c_10_p N_VSS_c_183_n 7.43603e-19
cc_34 N_VDD_c_11_p N_VSS_c_183_n 8.20353e-19
cc_35 N_VDD_c_16_p N_VSS_c_186_n 6.9475e-19
cc_36 N_VDD_c_21_p N_VSS_c_186_n 0.00161703f
cc_37 N_VDD_c_37_p N_VSS_c_186_n 9.10421e-19
cc_38 N_VDD_c_38_p N_VSS_c_186_n 3.48267e-19
cc_39 N_VDD_c_10_p N_VSS_c_190_n 4.06132e-19
cc_40 N_VDD_c_25_p N_VSS_c_190_n 0.00161703f
cc_41 N_VDD_c_11_p N_VSS_c_190_n 0.00146019f
cc_42 N_VDD_c_42_p N_VSS_c_190_n 3.48267e-19
cc_43 N_VDD_XI24.X0_PGD N_VSS_c_194_n 2.99706e-19
cc_44 N_VDD_c_37_p N_VSS_c_194_n 0.00524008f
cc_45 N_VDD_c_38_p N_VSS_c_194_n 9.58524e-19
cc_46 N_VDD_c_21_p N_VSS_c_197_n 0.00400652f
cc_47 N_VDD_c_13_p N_VSS_c_198_n 4.41003e-19
cc_48 N_VDD_c_30_p N_VSS_c_198_n 3.89161e-19
cc_49 N_VDD_c_2_p N_VSS_c_198_n 7.99831e-19
cc_50 N_VDD_c_16_p N_VSS_c_201_n 3.48267e-19
cc_51 N_VDD_c_21_p N_VSS_c_201_n 2.26455e-19
cc_52 N_VDD_c_37_p N_VSS_c_201_n 3.99794e-19
cc_53 N_VDD_c_38_p N_VSS_c_201_n 6.489e-19
cc_54 N_VDD_c_10_p N_VSS_c_205_n 3.82294e-19
cc_55 N_VDD_c_25_p N_VSS_c_205_n 2.26455e-19
cc_56 N_VDD_c_11_p N_VSS_c_205_n 9.55109e-19
cc_57 N_VDD_c_42_p N_VSS_c_205_n 6.46219e-19
cc_58 N_VDD_c_7_p N_VSS_c_209_n 0.00419405f
cc_59 N_VDD_c_13_p N_VSS_c_209_n 0.00325114f
cc_60 N_VDD_c_60_p N_VSS_c_209_n 0.0010705f
cc_61 N_VDD_c_13_p N_VSS_c_212_n 0.0102114f
cc_62 N_VDD_c_30_p N_VSS_c_212_n 0.00124944f
cc_63 N_VDD_c_5_p N_VSS_c_214_n 0.0097003f
cc_64 N_VDD_c_64_p N_VSS_c_215_n 0.00107633f
cc_65 N_VDD_c_65_p N_VSS_c_216_n 0.00833289f
cc_66 N_VDD_c_66_p N_VSS_c_216_n 6.51257e-19
cc_67 N_VDD_c_21_p N_VSS_c_216_n 0.00369311f
cc_68 N_VDD_c_68_p N_VSS_c_216_n 0.00146091f
cc_69 N_VDD_c_69_p N_VSS_c_220_n 0.00107845f
cc_70 N_VDD_c_5_p N_VSS_c_221_n 0.00143483f
cc_71 N_VDD_c_25_p N_VSS_c_221_n 0.00610315f
cc_72 N_VDD_c_72_p N_VSS_c_221_n 9.53204e-19
cc_73 N_VDD_c_10_p VSS 2.72347e-19
cc_74 N_VDD_c_11_p VSS 9.64592e-19
cc_75 N_VDD_c_13_p N_VSS_c_226_n 0.00109802f
cc_76 N_VDD_c_5_p N_VSS_c_227_n 0.00111918f
cc_77 N_VDD_c_21_p N_VSS_c_228_n 7.74609e-19
cc_78 N_VDD_c_78_p N_CI_c_285_n 3.43419e-19
cc_79 N_VDD_c_78_p N_CI_c_286_n 3.48267e-19
cc_80 N_VDD_c_5_p N_CI_c_286_n 3.21336e-19
cc_81 N_VDD_c_29_p N_CI_c_286_n 5.61123e-19
cc_82 N_VDD_c_30_p N_CI_c_286_n 0.00278407f
cc_83 N_VDD_c_16_p N_CI_c_290_n 7.63838e-19
cc_84 N_VDD_c_66_p N_CI_c_290_n 4.68699e-19
cc_85 N_VDD_XI24.X0_PGD N_A_c_332_n 3.96972e-19
cc_86 N_VDD_XI24.X0_PGD N_A_c_333_n 5.06189e-19
cc_87 N_VDD_c_6_p N_A_c_333_n 2.21087e-19
cc_88 N_VDD_c_21_p N_A_c_333_n 2.0692e-19
cc_89 N_VDD_c_11_p N_A_c_333_n 3.17218e-19
cc_90 N_VDD_c_38_p N_A_c_333_n 2.03128e-19
cc_91 N_VDD_c_6_p N_A_c_338_n 9.18655e-19
cc_92 N_VDD_c_11_p N_A_c_339_n 0.0068268f
cc_93 N_VDD_c_30_p N_A_c_340_n 0.00109781f
cc_94 N_VDD_c_30_p N_A_c_341_n 5.7233e-19
cc_95 N_VDD_c_6_p N_BI_c_401_n 3.43419e-19
cc_96 N_VDD_c_11_p N_BI_c_401_n 3.48267e-19
cc_97 N_VDD_c_6_p N_BI_c_403_n 3.48267e-19
cc_98 N_VDD_c_30_p N_BI_c_403_n 7.69656e-19
cc_99 N_VDD_c_25_p N_BI_c_403_n 3.21336e-19
cc_100 N_VDD_c_11_p N_BI_c_403_n 4.99861e-19
cc_101 N_VDD_XI24.X0_PGD N_AI_XI31.X0_PGD 3.10667e-19
cc_102 N_VDD_c_102_p N_AI_c_469_n 3.10667e-19
cc_103 N_VDD_c_103_p N_AI_c_470_n 3.43419e-19
cc_104 N_VDD_c_66_p N_AI_c_470_n 3.73302e-19
cc_105 N_VDD_c_103_p N_AI_c_472_n 3.48267e-19
cc_106 N_VDD_c_16_p N_AI_c_472_n 3.47482e-19
cc_107 N_VDD_c_66_p N_AI_c_472_n 5.23123e-19
cc_108 N_VDD_c_21_p N_AI_c_472_n 3.21336e-19
cc_109 N_VDD_c_37_p N_AI_c_476_n 0.00118673f
cc_110 N_VDD_XI26.X0_PGD N_B_XI25.X0_CG 0.00111782f
cc_111 N_VDD_XI25.X0_PGD N_B_c_515_n 4.01605e-19
cc_112 N_VDD_c_112_p N_B_c_516_n 0.00111782f
cc_113 N_VDD_c_11_p N_B_c_517_n 4.72333e-19
cc_114 N_C_c_116_n N_VSS_XI22.X0_PGD 4.20258e-19
cc_115 N_C_c_126_p N_VSS_c_230_n 2.76939e-19
cc_116 N_C_c_127_p N_VSS_c_183_n 7.31268e-19
cc_117 N_C_c_123_n N_VSS_c_183_n 0.00200258f
cc_118 N_C_c_129_p N_VSS_c_198_n 0.0041528f
cc_119 N_C_c_120_n N_VSS_c_209_n 4.01014e-19
cc_120 N_C_c_123_n N_VSS_c_209_n 2.67373e-19
cc_121 N_C_c_120_n N_VSS_c_214_n 0.00171716f
cc_122 N_C_c_123_n N_VSS_c_214_n 0.00318423f
cc_123 N_C_c_123_n N_VSS_c_221_n 0.00192963f
cc_124 N_C_c_123_n VSS 0.00167449f
cc_125 N_C_c_116_n N_CI_c_285_n 7.69306e-19
cc_126 N_C_c_123_n N_CI_c_286_n 7.42955e-19
cc_127 N_C_c_123_n N_CI_c_290_n 0.00148047f
cc_128 N_C_c_123_n N_A_c_333_n 3.38948e-19
cc_129 N_C_c_119_n N_A_c_338_n 8.20481e-19
cc_130 N_C_c_127_p N_A_c_338_n 0.00202163f
cc_131 N_C_c_123_n N_A_c_339_n 5.50651e-19
cc_132 N_C_c_143_p N_A_c_346_n 7.67297e-19
cc_133 N_C_c_119_n N_A_c_347_n 5.83331e-19
cc_134 N_C_c_127_p N_A_c_347_n 0.00118769f
cc_135 N_C_c_123_n N_A_c_347_n 4.69432e-19
cc_136 N_C_c_143_p N_A_c_347_n 0.00239654f
cc_137 N_C_c_148_p N_A_c_347_n 3.74525e-19
cc_138 N_C_c_123_n N_BI_c_403_n 2.74336e-19
cc_139 N_C_c_123_n N_BI_c_408_n 3.41448e-19
cc_140 N_C_c_143_p N_BI_c_409_n 4.45126e-19
cc_141 N_C_c_143_p N_BI_c_410_n 0.00127751f
cc_142 N_C_c_127_p N_B_c_517_n 0.00140507f
cc_143 N_C_c_123_n N_B_c_517_n 0.00214978f
cc_144 N_C_c_143_p N_B_c_517_n 9.13922e-19
cc_145 N_C_c_119_n N_Z_c_577_n 3.43419e-19
cc_146 N_C_c_157_p N_Z_c_577_n 3.43419e-19
cc_147 N_C_c_127_p N_Z_c_577_n 3.48267e-19
cc_148 N_C_c_159_p N_Z_c_577_n 3.48267e-19
cc_149 N_C_c_157_p N_Z_c_581_n 3.48267e-19
cc_150 N_C_c_127_p N_Z_c_581_n 6.09821e-19
cc_151 N_C_c_159_p N_Z_c_581_n 5.71987e-19
cc_152 N_VSS_c_177_n N_CI_c_285_n 3.43419e-19
cc_153 N_VSS_c_183_n N_CI_c_285_n 3.48267e-19
cc_154 N_VSS_c_242_p N_CI_c_297_n 3.43419e-19
cc_155 N_VSS_c_194_n N_CI_c_297_n 3.48267e-19
cc_156 N_VSS_c_177_n N_CI_c_286_n 3.48267e-19
cc_157 N_VSS_c_178_n N_CI_c_286_n 5.78167e-19
cc_158 N_VSS_c_183_n N_CI_c_286_n 0.00107566f
cc_159 N_VSS_c_209_n N_CI_c_286_n 6.53442e-19
cc_160 N_VSS_c_212_n N_CI_c_286_n 0.00285518f
cc_161 N_VSS_c_242_p N_CI_c_304_n 3.48267e-19
cc_162 N_VSS_c_194_n N_CI_c_304_n 0.00120696f
cc_163 N_VSS_c_186_n N_CI_c_290_n 0.00138401f
cc_164 N_VSS_c_194_n N_CI_c_290_n 2.05251e-19
cc_165 N_VSS_c_197_n N_CI_c_290_n 0.00334374f
cc_166 N_VSS_c_216_n N_CI_c_290_n 2.16087e-19
cc_167 N_VSS_c_216_n N_CI_c_310_n 0.00293637f
cc_168 N_VSS_XI21.X0_PGD N_A_c_332_n 3.96972e-19
cc_169 N_VSS_c_242_p N_A_c_333_n 4.13509e-19
cc_170 N_VSS_c_194_n N_A_c_333_n 7.30817e-19
cc_171 N_VSS_c_197_n N_A_c_333_n 2.62883e-19
cc_172 N_VSS_c_201_n N_A_c_340_n 2.09367e-19
cc_173 N_VSS_c_186_n N_A_c_341_n 2.04211e-19
cc_174 N_VSS_c_201_n N_A_c_341_n 4.89964e-19
cc_175 N_VSS_c_177_n N_BI_c_401_n 3.43419e-19
cc_176 N_VSS_c_183_n N_BI_c_401_n 3.48267e-19
cc_177 N_VSS_c_177_n N_BI_c_403_n 3.48267e-19
cc_178 N_VSS_c_183_n N_BI_c_403_n 0.00101872f
cc_179 N_VSS_c_221_n N_BI_c_403_n 2.19864e-19
cc_180 N_VSS_c_197_n N_BI_c_416_n 2.2551e-19
cc_181 N_VSS_XI23.X0_PGD N_AI_XI31.X0_PGD 2.79882e-19
cc_182 N_VSS_c_174_n N_AI_c_478_n 2.79882e-19
cc_183 N_VSS_c_242_p N_AI_c_470_n 3.43419e-19
cc_184 N_VSS_c_194_n N_AI_c_470_n 3.48267e-19
cc_185 N_VSS_c_242_p N_AI_c_472_n 3.48267e-19
cc_186 N_VSS_c_194_n N_AI_c_472_n 0.00173694f
cc_187 N_VSS_c_194_n N_AI_c_476_n 0.00177896f
cc_188 N_VSS_c_197_n N_AI_c_476_n 0.00605709f
cc_189 N_VSS_c_194_n N_AI_c_485_n 2.82216e-19
cc_190 N_VSS_c_186_n N_AI_c_486_n 0.00195338f
cc_191 N_VSS_c_197_n N_AI_c_486_n 0.00167789f
cc_192 N_VSS_XI23.X0_PGD N_B_c_515_n 4.01605e-19
cc_193 N_VSS_c_281_p N_B_c_522_n 6.24637e-19
cc_194 N_VSS_c_190_n B 2.2661e-19
cc_195 N_VSS_c_205_n B 2.39151e-19
cc_196 VSS N_B_c_517_n 2.35905e-19
cc_197 N_CI_c_290_n N_A_c_333_n 3.7003e-19
cc_198 N_CI_c_286_n N_BI_c_403_n 0.00144806f
cc_199 N_CI_c_313_p N_BI_c_418_n 5.10764e-19
cc_200 N_CI_c_304_n N_BI_c_408_n 6.46554e-19
cc_201 N_CI_c_290_n N_BI_c_408_n 8.14649e-19
cc_202 N_CI_c_313_p N_BI_c_409_n 0.0012701f
cc_203 N_CI_c_286_n N_AI_c_472_n 8.00553e-19
cc_204 N_CI_c_304_n N_AI_c_472_n 9.98055e-19
cc_205 N_CI_c_304_n N_AI_c_476_n 0.00117248f
cc_206 N_CI_c_290_n N_AI_c_476_n 0.00763297f
cc_207 N_CI_c_313_p N_AI_c_476_n 0.00313643f
cc_208 N_CI_c_322_p N_AI_c_476_n 0.00100316f
cc_209 N_CI_c_290_n N_AI_c_486_n 9.91646e-19
cc_210 N_CI_c_313_p N_B_c_526_n 7.08144e-19
cc_211 N_CI_c_297_n N_Z_c_584_n 3.43419e-19
cc_212 N_CI_c_326_p N_Z_c_584_n 3.43419e-19
cc_213 N_CI_c_304_n N_Z_c_584_n 3.48267e-19
cc_214 N_CI_c_328_p N_Z_c_584_n 3.48267e-19
cc_215 N_CI_c_326_p N_Z_c_581_n 3.48267e-19
cc_216 N_CI_c_304_n N_Z_c_581_n 6.09821e-19
cc_217 N_CI_c_328_p N_Z_c_581_n 5.71987e-19
cc_218 N_A_XI29.X0_PGD N_BI_XI29.X0_CG 9.65637e-19
cc_219 N_A_c_361_p N_BI_c_423_n 5.35095e-19
cc_220 N_A_c_333_n N_BI_c_403_n 3.00325e-19
cc_221 N_A_c_338_n N_BI_c_403_n 0.00110499f
cc_222 N_A_c_364_p N_BI_c_418_n 2.15082e-19
cc_223 N_A_XI29.X0_PGD N_BI_c_427_n 0.00133285f
cc_224 N_A_c_346_n N_BI_c_427_n 2.15082e-19
cc_225 N_A_c_338_n N_BI_c_408_n 0.00187419f
cc_226 N_A_c_333_n N_BI_c_416_n 0.00339867f
cc_227 N_A_c_338_n N_BI_c_431_n 3.69994e-19
cc_228 N_A_XI29.X0_PGD N_AI_XI31.X0_PGD 0.0173493f
cc_229 N_A_c_338_n N_AI_XI31.X0_PGD 0.001002f
cc_230 N_A_c_347_n N_AI_XI31.X0_PGD 7.67512e-19
cc_231 N_A_c_373_p N_AI_c_478_n 0.00199603f
cc_232 N_A_c_347_n N_AI_c_478_n 0.00128901f
cc_233 N_A_c_375_p N_AI_c_469_n 0.00201004f
cc_234 N_A_c_332_n N_AI_c_470_n 6.90199e-19
cc_235 N_A_c_333_n N_AI_c_472_n 5.84011e-19
cc_236 N_A_c_333_n N_AI_c_476_n 0.00127614f
cc_237 N_A_c_332_n N_B_c_515_n 0.00360349f
cc_238 N_A_c_333_n N_B_c_515_n 5.25071e-19
cc_239 N_A_c_340_n N_B_c_516_n 5.25071e-19
cc_240 N_A_c_341_n N_B_c_516_n 7.41063e-19
cc_241 N_A_c_333_n N_B_c_522_n 3.90215e-19
cc_242 N_A_XI29.X0_PGD N_B_c_532_n 9.65637e-19
cc_243 N_A_c_333_n B 6.34584e-19
cc_244 N_A_c_338_n B 4.3123e-19
cc_245 N_A_c_338_n N_B_c_535_n 4.01937e-19
cc_246 N_A_c_347_n N_B_c_535_n 3.79361e-19
cc_247 N_A_c_332_n N_B_c_537_n 7.73422e-19
cc_248 N_A_c_333_n N_B_c_537_n 5.77217e-19
cc_249 N_A_c_338_n N_B_c_537_n 6.37149e-19
cc_250 N_A_c_338_n N_B_c_540_n 3.37713e-19
cc_251 N_A_c_347_n N_B_c_540_n 2.21087e-19
cc_252 N_A_XI29.X0_PGD N_B_c_542_n 0.00133285f
cc_253 N_A_c_338_n N_B_c_517_n 0.00197838f
cc_254 N_A_c_347_n N_B_c_517_n 0.00180845f
cc_255 N_A_c_347_n N_Z_c_577_n 7.79328e-19
cc_256 N_A_XI29.X0_PGD N_Z_c_581_n 7.77706e-19
cc_257 N_A_c_338_n N_Z_c_581_n 0.00169143f
cc_258 N_A_c_347_n N_Z_c_581_n 0.0010247f
cc_259 N_BI_c_432_p N_AI_XI31.X0_PGD 9.65637e-19
cc_260 N_BI_c_433_p N_AI_XI31.X0_PGD 0.00133285f
cc_261 N_BI_c_416_n N_AI_c_472_n 6.07277e-19
cc_262 N_BI_c_433_p N_AI_c_476_n 2.15082e-19
cc_263 N_BI_c_408_n N_AI_c_476_n 0.00233431f
cc_264 N_BI_c_437_p N_AI_c_485_n 2.15082e-19
cc_265 N_BI_c_433_p N_AI_c_485_n 5.05931e-19
cc_266 N_BI_c_401_n N_B_c_515_n 6.90199e-19
cc_267 N_BI_c_403_n B 5.19468e-19
cc_268 N_BI_c_408_n B 2.66639e-19
cc_269 N_BI_c_437_p N_B_c_535_n 3.94971e-19
cc_270 N_BI_c_433_p N_B_c_535_n 4.03665e-19
cc_271 N_BI_c_408_n N_B_c_535_n 2.81186e-19
cc_272 N_BI_c_418_n N_B_c_526_n 0.00181951f
cc_273 N_BI_c_427_n N_B_c_526_n 4.56568e-19
cc_274 N_BI_c_437_p N_B_c_540_n 4.44913e-19
cc_275 N_BI_c_433_p N_B_c_540_n 0.00360065f
cc_276 N_BI_c_427_n N_B_c_540_n 0.00102603f
cc_277 N_BI_c_433_p N_B_c_542_n 7.16621e-19
cc_278 N_BI_c_427_n N_B_c_542_n 0.00243716f
cc_279 N_BI_c_403_n N_B_c_517_n 0.00150424f
cc_280 N_BI_c_418_n N_B_c_517_n 0.00163797f
cc_281 N_BI_c_408_n N_B_c_517_n 0.0161531f
cc_282 N_BI_c_409_n N_B_c_517_n 8.58649e-19
cc_283 N_BI_c_410_n N_B_c_517_n 6.57534e-19
cc_284 N_BI_c_408_n N_B_c_563_n 0.0022474f
cc_285 N_BI_c_458_p N_B_c_563_n 0.00206348f
cc_286 N_BI_c_410_n N_B_c_563_n 2.41136e-19
cc_287 N_BI_c_437_p N_B_c_566_n 3.09421e-19
cc_288 N_BI_c_431_n N_B_c_566_n 0.0022474f
cc_289 N_BI_c_409_n N_B_c_566_n 8.20948e-19
cc_290 N_BI_c_437_p N_Z_c_581_n 0.00157325f
cc_291 N_BI_c_418_n N_Z_c_581_n 0.00155051f
cc_292 N_BI_c_433_p N_Z_c_581_n 8.66889e-19
cc_293 N_BI_c_427_n N_Z_c_581_n 8.66889e-19
cc_294 N_BI_c_408_n N_Z_c_581_n 3.95297e-19
cc_295 N_AI_XI31.X0_PGD N_B_XI31.X0_CG 9.47088e-19
cc_296 N_AI_XI31.X0_PGD N_B_c_540_n 0.00340539f
cc_297 N_AI_XI31.X0_PGD N_Z_c_581_n 4.24987e-19
cc_298 N_B_c_535_n N_Z_c_581_n 0.00158441f
cc_299 N_B_c_526_n N_Z_c_581_n 0.00138952f
cc_300 N_B_c_542_n N_Z_c_581_n 8.66889e-19
cc_301 N_B_c_517_n N_Z_c_581_n 7.81804e-19
cc_302 N_B_c_563_n N_Z_c_581_n 0.00232585f
cc_303 N_B_c_566_n N_Z_c_581_n 0.00104129f
*
.ends
*
*
.subckt XNOR3_HPNW12 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XNOR3_N3
.ends
*
* File: G4_XOR2_N3.pex.netlist
* Created: Sun Apr 10 19:09:34 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G4_XOR2_N3_VSS 2 5 9 12 14 16 32 33 42 43 54 59 63 66 71 76 81 86 95
+ 100 113 115 116 117 122 123 128 138 140 145 146 147 150 Vss
c92 148 Vss 6.20041e-19
c93 147 Vss 3.75522e-19
c94 146 Vss 4.28045e-19
c95 145 Vss 0.00444873f
c96 140 Vss 0.00219072f
c97 138 Vss 0.00853623f
c98 128 Vss 0.00370986f
c99 123 Vss 8.46757e-19
c100 122 Vss 0.00174135f
c101 117 Vss 8.2479e-19
c102 116 Vss 0.00447709f
c103 115 Vss 0.00650684f
c104 113 Vss 0.00239513f
c105 100 Vss 0.00529998f
c106 95 Vss 0.00418654f
c107 86 Vss 2.86598e-19
c108 81 Vss 0.00160268f
c109 76 Vss 0.0010261f
c110 71 Vss 0.00123398f
c111 66 Vss 0.00174721f
c112 63 Vss 0.0101876f
c113 59 Vss 0.00691967f
c114 54 Vss 0.0100924f
c115 43 Vss 0.0342915f
c116 42 Vss 0.100071f
c117 33 Vss 0.0350852f
c118 32 Vss 0.0990727f
c119 14 Vss 0.00143493f
c120 9 Vss 0.384391f
c121 5 Vss 0.378692f
r122 145 150 0.326018
r123 144 145 5.50157
r124 140 144 0.655813
r125 139 148 0.494161
r126 138 150 0.326018
r127 138 139 13.0037
r128 134 148 0.128424
r129 129 147 0.494161
r130 128 148 0.494161
r131 128 129 7.46046
r132 124 147 0.128424
r133 122 147 0.494161
r134 122 123 4.37625
r135 118 146 0.0828784
r136 116 130 0.652036
r137 116 117 10.1279
r138 115 123 0.652036
r139 114 146 0.551426
r140 114 115 17.1716
r141 113 146 0.551426
r142 112 117 0.652036
r143 112 113 5.79332
r144 86 140 1.82344
r145 81 134 6.16843
r146 76 100 1.16709
r147 76 130 2.16729
r148 71 95 1.16709
r149 71 124 2.16729
r150 66 118 1.82344
r151 63 86 1.16709
r152 59 81 1.16709
r153 54 66 1.16709
r154 45 100 0.119107
r155 43 45 1.45875
r156 42 46 0.652036
r157 42 45 1.45875
r158 39 43 0.652036
r159 35 95 0.0476429
r160 33 35 1.45875
r161 32 36 0.652036
r162 32 35 1.45875
r163 29 33 0.652036
r164 16 63 0.123773
r165 14 59 0.123773
r166 12 59 0.123773
r167 9 46 5.1348
r168 9 39 5.1348
r169 5 36 5.1348
r170 5 29 5.1348
r171 2 54 0.123773
.ends

.subckt PM_G4_XOR2_N3_VDD 3 6 8 11 14 16 32 42 43 54 59 66 68 69 70 73 75 76 79
+ 81 85 89 91 93 98 99 100 103 109 114 123 Vss
c98 123 Vss 0.00813195f
c99 114 Vss 0.00444328f
c100 109 Vss 0.00562387f
c101 101 Vss 8.87755e-19
c102 100 Vss 2.39889e-19
c103 99 Vss 4.52364e-19
c104 98 Vss 0.0063791f
c105 93 Vss 0.00162315f
c106 91 Vss 0.0131786f
c107 89 Vss 0.00230903f
c108 85 Vss 7.1324e-19
c109 81 Vss 0.00459876f
c110 79 Vss 0.00140429f
c111 76 Vss 8.64616e-19
c112 75 Vss 0.00587269f
c113 73 Vss 0.00191373f
c114 70 Vss 8.68689e-19
c115 69 Vss 0.00224797f
c116 68 Vss 0.00279777f
c117 66 Vss 0.0108403f
c118 59 Vss 0.00695462f
c119 54 Vss 0.00822951f
c120 43 Vss 0.0351405f
c121 42 Vss 0.100972f
c122 33 Vss 0.0359366f
c123 32 Vss 0.100971f
c124 14 Vss 0.00143493f
c125 11 Vss 0.377105f
c126 3 Vss 0.384936f
r127 98 103 0.349767
r128 97 98 5.75164
r129 95 123 1.16709
r130 93 103 0.306046
r131 93 95 1.82344
r132 92 101 0.494161
r133 91 97 0.652036
r134 91 92 13.0037
r135 87 101 0.128424
r136 87 89 6.46018
r137 85 114 1.16709
r138 83 85 2.16729
r139 82 100 0.494161
r140 81 101 0.494161
r141 81 82 7.46046
r142 79 109 1.16709
r143 77 100 0.128424
r144 77 79 2.16729
r145 75 83 0.652036
r146 75 76 10.1279
r147 71 99 0.0828784
r148 71 73 1.82344
r149 69 100 0.494161
r150 69 70 4.37625
r151 68 76 0.652036
r152 67 99 0.551426
r153 67 68 5.50157
r154 66 99 0.551426
r155 65 70 0.652036
r156 65 66 17.4633
r157 63 123 0.05
r158 59 89 1.16709
r159 54 73 1.02121
r160 45 114 0.0476429
r161 43 45 1.45875
r162 42 46 0.652036
r163 42 45 1.45875
r164 39 43 0.652036
r165 35 109 0.119107
r166 33 35 1.45875
r167 32 36 0.652036
r168 32 35 1.45875
r169 29 33 0.652036
r170 16 63 0.123773
r171 14 59 0.123773
r172 11 46 5.1348
r173 11 39 5.1348
r174 8 59 0.123773
r175 6 54 0.123773
r176 3 36 5.1348
r177 3 29 5.1348
.ends

.subckt PM_G4_XOR2_N3_A 2 4 7 10 21 24 28 48 51 54 57 62 67 72 77 85 Vss
c54 85 Vss 8.24403e-19
c55 77 Vss 0.00191043f
c56 72 Vss 0.00680655f
c57 67 Vss 0.00366581f
c58 62 Vss 0.00280314f
c59 57 Vss 0.00457389f
c60 51 Vss 0.00108099f
c61 48 Vss 0.128068f
c62 43 Vss 0.0296639f
c63 28 Vss 0.152693f
c64 24 Vss 8.47557e-20
c65 21 Vss 0.173351f
c66 18 Vss 0.180502f
c67 16 Vss 0.0247918f
c68 10 Vss 0.176342f
c69 7 Vss 0.432086f
c70 4 Vss 0.193054f
r71 81 85 0.653045
r72 62 77 1.16709
r73 62 85 4.9014
r74 57 72 1.16709
r75 57 81 10.8364
r76 51 67 1.16709
r77 51 54 0.0833571
r78 47 72 0.0238214
r79 47 48 2.334
r80 44 47 2.20433
r81 39 77 0.50025
r82 33 48 0.00605528
r83 31 44 0.00605528
r84 29 43 0.494161
r85 28 30 0.652036
r86 28 29 4.84305
r87 25 43 0.128424
r88 24 67 0.0476429
r89 22 24 0.326018
r90 22 24 0.1167
r91 21 43 0.494161
r92 21 24 6.7686
r93 18 67 0.357321
r94 16 24 0.326018
r95 16 18 0.40845
r96 10 39 4.668
r97 7 33 5.1348
r98 7 31 5.1348
r99 7 30 5.1348
r100 4 25 5.1348
r101 2 18 4.72635
.ends

.subckt PM_G4_XOR2_N3_NET1 2 4 7 10 31 35 41 44 49 58 76 Vss
c34 76 Vss 3.97901e-19
c35 58 Vss 0.0058132f
c36 49 Vss 0.00651255f
c37 44 Vss 0.00236298f
c38 41 Vss 0.00514975f
c39 35 Vss 0.103147f
c40 31 Vss 0.12549f
c41 10 Vss 0.269166f
c42 7 Vss 0.499657f
c43 4 Vss 0.00143493f
r44 72 76 0.655813
r45 49 58 1.16709
r46 49 76 12.1076
r47 44 72 3.62604
r48 41 44 1.16709
r49 33 35 1.70187
r50 30 58 0.142929
r51 30 31 2.20433
r52 27 30 2.334
r53 25 35 0.17282
r54 24 31 0.00605528
r55 21 33 0.17282
r56 18 27 0.00605528
r57 10 21 7.64385
r58 7 25 7.29375
r59 7 24 5.1348
r60 7 18 5.1348
r61 4 41 0.123773
r62 2 41 0.123773
.ends

.subckt PM_G4_XOR2_N3_NET2 2 4 6 9 21 22 33 39 42 47 56 74 Vss
c42 74 Vss 3.21991e-19
c43 56 Vss 0.00502059f
c44 47 Vss 0.00781175f
c45 42 Vss 0.00242715f
c46 39 Vss 0.00509494f
c47 33 Vss 0.12909f
c48 22 Vss 0.0345713f
c49 21 Vss 0.177367f
c50 9 Vss 0.573605f
c51 6 Vss 0.188648f
c52 4 Vss 0.00143493f
r53 70 74 0.660011
r54 47 56 1.16709
r55 47 74 11.3611
r56 42 70 3.29261
r57 39 42 1.16709
r58 32 56 0.0238214
r59 32 33 2.26917
r60 29 32 2.26917
r61 26 33 0.00605528
r62 24 29 0.00605528
r63 21 23 0.652036
r64 21 22 4.84305
r65 18 22 0.652036
r66 9 26 5.1348
r67 9 24 5.1348
r68 9 23 10.0362
r69 6 18 5.1348
r70 4 39 0.123773
r71 2 39 0.123773
.ends

.subckt PM_G4_XOR2_N3_B 2 4 7 10 19 20 28 31 35 45 51 54 Vss
c31 54 Vss 0.0283542f
c32 51 Vss 0.00177471f
c33 45 Vss 0.13328f
c34 35 Vss 0.154928f
c35 31 Vss 2.04877e-19
c36 28 Vss 0.117534f
c37 20 Vss 0.0348422f
c38 19 Vss 0.173065f
c39 10 Vss 0.264298f
c40 7 Vss 0.440555f
c41 4 Vss 0.189408f
c42 2 Vss 0.201403f
r43 51 54 1.16709
r44 43 45 4.53833
r45 38 45 0.00605528
r46 35 47 1.87725
r47 33 47 0.527901
r48 32 43 0.00605528
r49 31 54 0.181909
r50 29 54 0.494161
r51 29 31 0.1167
r52 28 47 0.333556
r53 28 31 4.72635
r54 23 54 0.128424
r55 23 54 0.40845
r56 22 54 0.181909
r57 20 22 6.7686
r58 19 54 0.494161
r59 19 22 0.1167
r60 16 20 0.652036
r61 10 35 7.5855
r62 7 38 5.1348
r63 7 33 5.42655
r64 7 32 5.1348
r65 4 54 5.0181
r66 2 16 5.42655
.ends

.subckt PM_G4_XOR2_N3_Z 2 4 6 8 23 27 30 33 Vss
c29 30 Vss 0.00322833f
c30 27 Vss 0.00675283f
c31 23 Vss 0.00497092f
c32 8 Vss 0.00143493f
c33 6 Vss 0.00143493f
r34 33 35 4.95975
r35 30 33 6.71025
r36 27 35 1.16709
r37 23 30 1.16709
r38 8 27 0.123773
r39 6 23 0.123773
r40 4 27 0.123773
r41 2 23 0.123773
.ends

.subckt G4_XOR2_N3  VSS VDD A B Z
*
* Z	Z
* B	B
* A	A
* VDD	VDD
* VSS	VSS
XI20.X0 N_NET1_XI20.X0_D N_VDD_XI20.X0_PGD N_B_XI20.X0_CG N_VDD_XI20.X0_PGD
+ N_VSS_XI20.X0_S TIGFET_HPNW12
XI18.X0 N_NET2_XI18.X0_D N_VSS_XI18.X0_PGD N_A_XI18.X0_CG N_VSS_XI18.X0_PGD
+ N_VDD_XI18.X0_S TIGFET_HPNW12
XI22.X0 N_NET1_XI22.X0_D N_VSS_XI22.X0_PGD N_B_XI22.X0_CG N_VSS_XI22.X0_PGD
+ N_VDD_XI22.X0_S TIGFET_HPNW12
XI16.X0 N_NET2_XI16.X0_D N_VDD_XI16.X0_PGD N_A_XI16.X0_CG N_VDD_XI16.X0_PGD
+ N_VSS_XI16.X0_S TIGFET_HPNW12
XI21.X0 N_Z_XI21.X0_D N_B_XI21.X0_PGD N_NET2_XI21.X0_CG N_B_XI21.X0_PGD
+ N_VDD_XI21.X0_S TIGFET_HPNW12
XI19.X0 N_Z_XI19.X0_D N_A_XI19.X0_PGD N_B_XI19.X0_CG N_A_XI19.X0_PGD
+ N_VSS_XI19.X0_S TIGFET_HPNW12
XI23.X0 N_Z_XI23.X0_D N_NET1_XI23.X0_PGD N_A_XI23.X0_CG N_NET1_XI23.X0_PGD
+ N_VDD_XI23.X0_S TIGFET_HPNW12
XI17.X0 N_Z_XI17.X0_D N_NET2_XI17.X0_PGD N_NET1_XI17.X0_CG N_NET2_XI17.X0_PGD
+ N_VSS_XI17.X0_S TIGFET_HPNW12
*
x_PM_G4_XOR2_N3_VSS N_VSS_XI20.X0_S N_VSS_XI18.X0_PGD N_VSS_XI22.X0_PGD
+ N_VSS_XI16.X0_S N_VSS_XI19.X0_S N_VSS_XI17.X0_S N_VSS_c_5_p N_VSS_c_22_p
+ N_VSS_c_38_p N_VSS_c_4_p N_VSS_c_7_p N_VSS_c_6_p N_VSS_c_85_p N_VSS_c_8_p
+ N_VSS_c_13_p N_VSS_c_29_p N_VSS_c_36_p N_VSS_c_87_p N_VSS_c_14_p N_VSS_c_30_p
+ N_VSS_c_9_p N_VSS_c_10_p N_VSS_c_18_p N_VSS_c_19_p N_VSS_c_25_p N_VSS_c_28_p
+ N_VSS_c_26_p N_VSS_c_55_p N_VSS_c_41_p N_VSS_c_57_p N_VSS_c_11_p N_VSS_c_27_p
+ VSS Vss PM_G4_XOR2_N3_VSS
x_PM_G4_XOR2_N3_VDD N_VDD_XI20.X0_PGD N_VDD_XI18.X0_S N_VDD_XI22.X0_S
+ N_VDD_XI16.X0_PGD N_VDD_XI21.X0_S N_VDD_XI23.X0_S N_VDD_c_96_n N_VDD_c_144_p
+ N_VDD_c_97_n N_VDD_c_167_p N_VDD_c_98_n N_VDD_c_99_n N_VDD_c_104_n
+ N_VDD_c_108_n N_VDD_c_111_n N_VDD_c_112_n N_VDD_c_113_n N_VDD_c_120_n
+ N_VDD_c_121_n N_VDD_c_123_n N_VDD_c_127_n N_VDD_c_130_n N_VDD_c_148_p
+ N_VDD_c_133_n N_VDD_c_155_p N_VDD_c_134_n N_VDD_c_135_n VDD N_VDD_c_136_n
+ N_VDD_c_138_n N_VDD_c_185_p Vss PM_G4_XOR2_N3_VDD
x_PM_G4_XOR2_N3_A N_A_XI18.X0_CG N_A_XI16.X0_CG N_A_XI19.X0_PGD N_A_XI23.X0_CG
+ N_A_c_191_n N_A_c_193_n N_A_c_194_n N_A_c_208_n N_A_c_195_n A N_A_c_196_n
+ N_A_c_201_n N_A_c_202_n N_A_c_215_n N_A_c_219_p N_A_c_203_n Vss
+ PM_G4_XOR2_N3_A
x_PM_G4_XOR2_N3_NET1 N_NET1_XI20.X0_D N_NET1_XI22.X0_D N_NET1_XI23.X0_PGD
+ N_NET1_XI17.X0_CG N_NET1_c_250_n N_NET1_c_270_p N_NET1_c_245_n N_NET1_c_246_n
+ N_NET1_c_247_n N_NET1_c_259_n N_NET1_c_248_n Vss PM_G4_XOR2_N3_NET1
x_PM_G4_XOR2_N3_NET2 N_NET2_XI18.X0_D N_NET2_XI16.X0_D N_NET2_XI21.X0_CG
+ N_NET2_XI17.X0_PGD N_NET2_c_300_n N_NET2_c_315_p N_NET2_c_301_n N_NET2_c_279_n
+ N_NET2_c_281_n N_NET2_c_284_n N_NET2_c_306_n N_NET2_c_288_n Vss
+ PM_G4_XOR2_N3_NET2
x_PM_G4_XOR2_N3_B N_B_XI20.X0_CG N_B_XI22.X0_CG N_B_XI21.X0_PGD N_B_XI19.X0_CG
+ N_B_c_323_n N_B_c_338_n N_B_c_325_n N_B_c_326_n N_B_c_340_n N_B_c_327_n B
+ N_B_c_335_n Vss PM_G4_XOR2_N3_B
x_PM_G4_XOR2_N3_Z N_Z_XI21.X0_D N_Z_XI19.X0_D N_Z_XI23.X0_D N_Z_XI17.X0_D
+ N_Z_c_361_n N_Z_c_352_n N_Z_c_356_n Z Vss PM_G4_XOR2_N3_Z
cc_1 N_VSS_XI18.X0_PGD N_VDD_XI20.X0_PGD 3.18967e-19
cc_2 N_VSS_XI22.X0_PGD N_VDD_XI20.X0_PGD 0.00194647f
cc_3 N_VSS_XI18.X0_PGD N_VDD_XI16.X0_PGD 0.00196596f
cc_4 N_VSS_c_4_p N_VDD_c_96_n 0.00194647f
cc_5 N_VSS_c_5_p N_VDD_c_97_n 0.00196596f
cc_6 N_VSS_c_6_p N_VDD_c_98_n 3.76525e-19
cc_7 N_VSS_c_7_p N_VDD_c_99_n 9.5668e-19
cc_8 N_VSS_c_8_p N_VDD_c_99_n 0.00165395f
cc_9 N_VSS_c_9_p N_VDD_c_99_n 0.00452338f
cc_10 N_VSS_c_10_p N_VDD_c_99_n 0.00889981f
cc_11 N_VSS_c_11_p N_VDD_c_99_n 9.16632e-19
cc_12 N_VSS_XI18.X0_PGD N_VDD_c_104_n 3.80615e-19
cc_13 N_VSS_c_13_p N_VDD_c_104_n 4.35319e-19
cc_14 N_VSS_c_14_p N_VDD_c_104_n 3.66936e-19
cc_15 N_VSS_c_10_p N_VDD_c_104_n 0.0039632f
cc_16 N_VSS_c_7_p N_VDD_c_108_n 2.57623e-19
cc_17 N_VSS_c_8_p N_VDD_c_108_n 3.02798e-19
cc_18 N_VSS_c_18_p N_VDD_c_108_n 0.00357068f
cc_19 N_VSS_c_19_p N_VDD_c_111_n 0.00106367f
cc_20 N_VSS_c_8_p N_VDD_c_112_n 4.43088e-19
cc_21 N_VSS_c_5_p N_VDD_c_113_n 3.89167e-19
cc_22 N_VSS_c_22_p N_VDD_c_113_n 3.89167e-19
cc_23 N_VSS_c_13_p N_VDD_c_113_n 0.00161703f
cc_24 N_VSS_c_14_p N_VDD_c_113_n 2.26455e-19
cc_25 N_VSS_c_25_p N_VDD_c_113_n 0.00348402f
cc_26 N_VSS_c_26_p N_VDD_c_113_n 0.00600907f
cc_27 N_VSS_c_27_p N_VDD_c_113_n 7.74609e-19
cc_28 N_VSS_c_28_p N_VDD_c_120_n 0.00107963f
cc_29 N_VSS_c_29_p N_VDD_c_121_n 9.20609e-19
cc_30 N_VSS_c_30_p N_VDD_c_121_n 3.82294e-19
cc_31 N_VSS_c_4_p N_VDD_c_123_n 3.76472e-19
cc_32 N_VSS_c_29_p N_VDD_c_123_n 0.00141228f
cc_33 N_VSS_c_30_p N_VDD_c_123_n 0.00112249f
cc_34 N_VSS_c_18_p N_VDD_c_123_n 0.00616046f
cc_35 N_VSS_c_13_p N_VDD_c_127_n 9.25616e-19
cc_36 N_VSS_c_36_p N_VDD_c_127_n 8.475e-19
cc_37 N_VSS_c_14_p N_VDD_c_127_n 3.99794e-19
cc_38 N_VSS_c_38_p N_VDD_c_130_n 2.88732e-19
cc_39 N_VSS_c_29_p N_VDD_c_130_n 0.00232715f
cc_40 N_VSS_c_30_p N_VDD_c_130_n 9.55109e-19
cc_41 N_VSS_c_41_p N_VDD_c_133_n 9.21122e-19
cc_42 N_VSS_c_10_p N_VDD_c_134_n 0.0010705f
cc_43 N_VSS_c_18_p N_VDD_c_135_n 9.68246e-19
cc_44 N_VSS_c_29_p N_VDD_c_136_n 3.48267e-19
cc_45 N_VSS_c_30_p N_VDD_c_136_n 8.00903e-19
cc_46 N_VSS_c_13_p N_VDD_c_138_n 3.48267e-19
cc_47 N_VSS_c_14_p N_VDD_c_138_n 6.489e-19
cc_48 N_VSS_XI18.X0_PGD N_A_c_191_n 4.09718e-19
cc_49 N_VSS_XI22.X0_PGD N_A_c_191_n 2.49973e-19
cc_50 N_VSS_c_14_p N_A_c_193_n 5.35095e-19
cc_51 N_VSS_XI22.X0_PGD N_A_c_194_n 2.49973e-19
cc_52 N_VSS_c_14_p N_A_c_195_n 2.15082e-19
cc_53 N_VSS_c_36_p N_A_c_196_n 0.00705874f
cc_54 N_VSS_c_10_p N_A_c_196_n 9.14669e-19
cc_55 N_VSS_c_55_p N_A_c_196_n 0.00173435f
cc_56 N_VSS_c_41_p N_A_c_196_n 3.96468e-19
cc_57 N_VSS_c_57_p N_A_c_196_n 4.40676e-19
cc_58 N_VSS_c_55_p N_A_c_201_n 6.19395e-19
cc_59 N_VSS_c_13_p N_A_c_202_n 2.15082e-19
cc_60 N_VSS_c_55_p N_A_c_203_n 4.24683e-19
cc_61 N_VSS_c_7_p N_NET1_c_245_n 3.43419e-19
cc_62 N_VSS_c_8_p N_NET1_c_246_n 0.00115894f
cc_63 N_VSS_c_29_p N_NET1_c_247_n 0.00149535f
cc_64 N_VSS_c_9_p N_NET1_c_248_n 7.76947e-19
cc_65 N_VSS_c_18_p N_NET1_c_248_n 6.52479e-19
cc_66 N_VSS_c_6_p N_NET2_c_279_n 3.43419e-19
cc_67 N_VSS_c_36_p N_NET2_c_279_n 3.48267e-19
cc_68 N_VSS_c_6_p N_NET2_c_281_n 3.48267e-19
cc_69 N_VSS_c_36_p N_NET2_c_281_n 0.00192385f
cc_70 N_VSS_c_10_p N_NET2_c_281_n 8.02212e-19
cc_71 N_VSS_c_36_p N_NET2_c_284_n 0.00186158f
cc_72 N_VSS_c_26_p N_NET2_c_284_n 0.00117864f
cc_73 N_VSS_c_55_p N_NET2_c_284_n 0.00504587f
cc_74 N_VSS_c_57_p N_NET2_c_284_n 0.00115623f
cc_75 N_VSS_c_13_p N_NET2_c_288_n 5.67902e-19
cc_76 N_VSS_c_26_p N_NET2_c_288_n 4.84133e-19
cc_77 N_VSS_c_30_p N_B_XI22.X0_CG 0.00322194f
cc_78 N_VSS_XI22.X0_PGD N_B_XI21.X0_PGD 0.00189584f
cc_79 N_VSS_XI18.X0_PGD N_B_c_323_n 2.60477e-19
cc_80 N_VSS_XI22.X0_PGD N_B_c_323_n 4.09718e-19
cc_81 N_VSS_XI22.X0_PGD N_B_c_325_n 4.09718e-19
cc_82 N_VSS_c_30_p N_B_c_326_n 2.76939e-19
cc_83 N_VSS_c_38_p N_B_c_327_n 0.00167898f
cc_84 N_VSS_c_6_p N_Z_c_352_n 3.43419e-19
cc_85 N_VSS_c_85_p N_Z_c_352_n 3.43419e-19
cc_86 N_VSS_c_36_p N_Z_c_352_n 3.48267e-19
cc_87 N_VSS_c_87_p N_Z_c_352_n 3.48267e-19
cc_88 N_VSS_c_6_p N_Z_c_356_n 3.48267e-19
cc_89 N_VSS_c_85_p N_Z_c_356_n 3.48267e-19
cc_90 N_VSS_c_36_p N_Z_c_356_n 4.84964e-19
cc_91 N_VSS_c_87_p N_Z_c_356_n 5.71987e-19
cc_92 N_VSS_c_55_p N_Z_c_356_n 3.20264e-19
cc_93 N_VDD_XI16.X0_PGD N_A_XI19.X0_PGD 0.00169921f
cc_94 N_VDD_XI20.X0_PGD N_A_c_191_n 2.49973e-19
cc_95 N_VDD_XI16.X0_PGD N_A_c_191_n 4.09718e-19
cc_96 N_VDD_XI16.X0_PGD N_A_c_194_n 4.09718e-19
cc_97 N_VDD_c_144_p N_A_c_208_n 0.00169921f
cc_98 N_VDD_c_99_n N_A_c_195_n 5.04211e-19
cc_99 N_VDD_c_127_n N_A_c_196_n 5.50187e-19
cc_100 N_VDD_c_138_n N_A_c_196_n 3.5189e-19
cc_101 N_VDD_c_148_p N_A_c_201_n 5.4427e-19
cc_102 N_VDD_c_99_n N_A_c_202_n 6.25289e-19
cc_103 N_VDD_c_136_n N_A_c_202_n 2.53697e-19
cc_104 N_VDD_c_127_n N_A_c_215_n 4.08069e-19
cc_105 N_VDD_c_138_n N_A_c_215_n 6.61916e-19
cc_106 N_VDD_c_148_p N_A_c_203_n 7.25922e-19
cc_107 N_VDD_c_148_p N_NET1_c_250_n 8.20153e-19
cc_108 N_VDD_c_155_p N_NET1_c_250_n 4.09731e-19
cc_109 N_VDD_c_98_n N_NET1_c_245_n 3.43419e-19
cc_110 N_VDD_c_98_n N_NET1_c_246_n 3.48267e-19
cc_111 N_VDD_c_123_n N_NET1_c_246_n 2.9283e-19
cc_112 N_VDD_c_130_n N_NET1_c_246_n 0.00152282f
cc_113 N_VDD_c_130_n N_NET1_c_247_n 0.00160739f
cc_114 N_VDD_c_148_p N_NET1_c_247_n 0.00374811f
cc_115 N_VDD_c_155_p N_NET1_c_247_n 8.18723e-19
cc_116 N_VDD_c_130_n N_NET1_c_259_n 2.78343e-19
cc_117 N_VDD_c_148_p N_NET1_c_259_n 2.37583e-19
cc_118 N_VDD_c_155_p N_NET1_c_259_n 3.70842e-19
cc_119 N_VDD_c_121_n N_NET1_c_248_n 2.88872e-19
cc_120 N_VDD_c_167_p N_NET2_c_279_n 3.67949e-19
cc_121 N_VDD_c_112_n N_NET2_c_279_n 3.72199e-19
cc_122 N_VDD_c_167_p N_NET2_c_281_n 3.9802e-19
cc_123 N_VDD_c_112_n N_NET2_c_281_n 5.226e-19
cc_124 N_VDD_c_113_n N_NET2_c_281_n 3.21336e-19
cc_125 N_VDD_c_127_n N_NET2_c_284_n 3.20822e-19
cc_126 N_VDD_c_99_n N_B_XI20.X0_CG 3.86879e-19
cc_127 N_VDD_c_136_n N_B_XI20.X0_CG 0.00180351f
cc_128 N_VDD_XI20.X0_PGD N_B_c_323_n 4.09718e-19
cc_129 N_VDD_XI16.X0_PGD N_B_c_323_n 2.60477e-19
cc_130 N_VDD_XI16.X0_PGD N_B_c_325_n 2.60477e-19
cc_131 N_VDD_c_130_n N_B_c_327_n 3.02511e-19
cc_132 N_VDD_c_148_p N_B_c_327_n 9.69761e-19
cc_133 N_VDD_c_138_n N_B_c_335_n 4.47793e-19
cc_134 N_VDD_c_98_n N_Z_c_361_n 3.43419e-19
cc_135 N_VDD_c_130_n N_Z_c_361_n 3.48267e-19
cc_136 N_VDD_c_148_p N_Z_c_361_n 2.57623e-19
cc_137 N_VDD_c_133_n N_Z_c_361_n 3.72199e-19
cc_138 N_VDD_c_185_p N_Z_c_361_n 3.43419e-19
cc_139 N_VDD_c_98_n N_Z_c_356_n 3.48267e-19
cc_140 N_VDD_c_130_n N_Z_c_356_n 7.9714e-19
cc_141 N_VDD_c_148_p N_Z_c_356_n 4.72042e-19
cc_142 N_VDD_c_133_n N_Z_c_356_n 8.30519e-19
cc_143 N_VDD_c_185_p N_Z_c_356_n 3.48267e-19
cc_144 N_A_XI23.X0_CG N_NET1_XI23.X0_PGD 9.16948e-19
cc_145 N_A_c_219_p N_NET1_XI23.X0_PGD 9.43732e-19
cc_146 N_A_c_201_n N_NET1_c_247_n 0.00175052f
cc_147 N_A_c_203_n N_NET1_c_247_n 5.83558e-19
cc_148 N_A_XI23.X0_CG N_NET1_c_259_n 0.00320789f
cc_149 N_A_c_219_p N_NET1_c_259_n 4.20251e-19
cc_150 N_A_XI23.X0_CG N_NET2_XI21.X0_CG 2.29068e-19
cc_151 N_A_XI19.X0_PGD N_NET2_XI17.X0_PGD 0.00174694f
cc_152 N_A_c_194_n N_NET2_XI17.X0_PGD 3.14428e-19
cc_153 N_A_c_219_p N_NET2_XI17.X0_PGD 3.71891e-19
cc_154 N_A_XI19.X0_PGD N_NET2_c_300_n 4.64512e-19
cc_155 N_A_c_208_n N_NET2_c_301_n 0.00174694f
cc_156 N_A_c_191_n N_NET2_c_279_n 6.03094e-19
cc_157 N_A_c_196_n N_NET2_c_284_n 0.002281f
cc_158 N_A_c_201_n N_NET2_c_284_n 9.32615e-19
cc_159 N_A_c_215_n N_NET2_c_284_n 3.44698e-19
cc_160 N_A_c_196_n N_NET2_c_306_n 3.44698e-19
cc_161 N_A_c_215_n N_NET2_c_306_n 6.78604e-19
cc_162 N_A_c_194_n N_B_XI19.X0_CG 0.003858f
cc_163 N_A_c_191_n N_B_c_323_n 0.00635057f
cc_164 N_A_c_202_n N_B_c_338_n 9.89912e-19
cc_165 N_A_c_194_n N_B_c_325_n 0.00470625f
cc_166 N_A_c_194_n N_B_c_340_n 0.00225174f
cc_167 N_A_c_191_n N_B_c_335_n 0.00106939f
cc_168 N_A_c_196_n N_Z_c_356_n 0.00384185f
cc_169 N_A_c_201_n N_Z_c_356_n 0.00366674f
cc_170 N_A_c_219_p N_Z_c_356_n 9.50702e-19
cc_171 N_NET1_XI23.X0_PGD N_NET2_XI21.X0_CG 2.3921e-19
cc_172 N_NET1_c_270_p N_NET2_XI17.X0_PGD 0.00794356f
cc_173 N_NET1_XI23.X0_PGD N_NET2_c_300_n 0.00388625f
cc_174 N_NET1_c_245_n N_NET2_c_279_n 2.80316e-19
cc_175 N_NET1_XI23.X0_PGD N_B_XI21.X0_PGD 0.00215617f
cc_176 N_NET1_XI17.X0_CG N_B_XI19.X0_CG 2.58346e-19
cc_177 N_NET1_c_245_n N_B_c_323_n 5.56563e-19
cc_178 N_NET1_c_270_p N_B_c_340_n 2.58346e-19
cc_179 N_NET1_c_250_n N_B_c_327_n 0.00193019f
cc_180 N_NET1_c_247_n N_Z_c_356_n 2.27374e-19
cc_181 N_NET2_XI21.X0_CG N_B_XI21.X0_PGD 0.00204226f
cc_182 N_NET2_c_300_n N_B_XI21.X0_PGD 0.00163867f
cc_183 N_NET2_XI17.X0_PGD N_B_c_340_n 0.00351134f
cc_184 N_NET2_c_315_p N_B_c_340_n 0.00405072f
cc_185 N_NET2_c_300_n N_Z_c_361_n 7.50005e-19
cc_186 N_NET2_c_300_n N_Z_c_352_n 2.48148e-19
cc_187 N_NET2_XI17.X0_PGD N_Z_c_356_n 0.00113722f
cc_188 N_NET2_c_300_n N_Z_c_356_n 2.5304e-19
cc_189 N_NET2_c_284_n N_Z_c_356_n 3.45637e-19
cc_190 N_B_c_340_n N_Z_c_356_n 0.00106974f
*
.ends
*
*
.subckt XOR2_HPNW12 A B Y VDD VSS
xgate (VSS VDD A B Y) G4_XOR2_N3
.ends
*
* File: G5_XOR3_N3.pex.netlist
* Created: Fri Apr  1 15:48:12 2022
* Program "Calibre xRC"
* Version "v2021.2_37.20"
*
.subckt PM_G5_XOR3_N3_VDD 2 5 9 12 14 17 34 35 44 45 54 55 65 69 74 77 79 80 81
+ 84 86 90 93 96 98 102 104 108 112 114 116 118 119 125 134 139 Vss
c113 139 Vss 0.00510833f
c114 134 Vss 0.00495479f
c115 125 Vss 0.00566756f
c116 119 Vss 2.39889e-19
c117 118 Vss 4.92173e-19
c118 117 Vss 5.50975e-19
c119 114 Vss 4.52364e-19
c120 112 Vss 0.00180866f
c121 108 Vss 0.00116218f
c122 104 Vss 0.00632073f
c123 102 Vss 0.0010418f
c124 98 Vss 0.00598007f
c125 96 Vss 0.00126332f
c126 93 Vss 0.00323042f
c127 90 Vss 0.00584753f
c128 86 Vss 0.00654417f
c129 84 Vss 0.00154142f
c130 81 Vss 8.68392e-19
c131 80 Vss 0.00938293f
c132 79 Vss 0.0122224f
c133 77 Vss 0.00304889f
c134 74 Vss 0.00820121f
c135 69 Vss 0.00836757f
c136 65 Vss 0.00811483f
c137 55 Vss 0.0356247f
c138 54 Vss 0.10084f
c139 45 Vss 0.0356281f
c140 44 Vss 0.101312f
c141 35 Vss 0.0346562f
c142 34 Vss 0.0991017f
c143 17 Vss 0.378774f
c144 9 Vss 0.379342f
c145 5 Vss 0.383323f
r146 110 112 6.16843
r147 108 139 1.16709
r148 106 108 2.16729
r149 105 119 0.494161
r150 104 110 0.652036
r151 104 105 7.46046
r152 102 134 1.16709
r153 100 119 0.128424
r154 100 102 2.16729
r155 99 118 0.494161
r156 98 106 0.652036
r157 98 99 10.3363
r158 94 117 0.0828784
r159 94 96 2.00578
r160 93 118 0.128424
r161 92 117 0.551426
r162 92 93 5.50157
r163 90 125 1.16709
r164 88 117 0.551426
r165 88 90 7.66886
r166 87 116 0.326018
r167 86 118 0.494161
r168 86 87 10.1279
r169 82 114 0.0828784
r170 82 84 1.82344
r171 80 119 0.494161
r172 80 81 15.8795
r173 79 116 0.326018
r174 78 114 0.551426
r175 78 79 18.3386
r176 77 114 0.551426
r177 76 81 0.652036
r178 76 77 5.50157
r179 74 112 1.16709
r180 69 96 1.16709
r181 65 84 1.16709
r182 57 139 0.0476429
r183 55 57 1.45875
r184 54 58 0.652036
r185 54 57 1.45875
r186 51 55 0.652036
r187 47 134 0.0476429
r188 45 47 1.45875
r189 44 48 0.652036
r190 44 47 1.45875
r191 41 45 0.652036
r192 37 125 0.238214
r193 35 37 1.45875
r194 34 38 0.652036
r195 34 37 1.45875
r196 31 35 0.652036
r197 17 58 5.1348
r198 17 51 5.1348
r199 14 74 0.123773
r200 12 69 0.123773
r201 9 48 5.1348
r202 9 41 5.1348
r203 5 38 5.1348
r204 5 31 5.1348
r205 2 65 0.123773
.ends

.subckt PM_G5_XOR3_N3_C 2 4 6 8 17 20 23 32 37 40 44 47 52 57 84 92 98 Vss
c49 98 Vss 3.22849e-19
c50 92 Vss 0.00543331f
c51 84 Vss 0.00847968f
c52 57 Vss 0.004971f
c53 52 Vss 7.31044e-19
c54 47 Vss 9.97921e-19
c55 40 Vss 0.00163759f
c56 37 Vss 0.0082356f
c57 32 Vss 0.00958317f
c58 23 Vss 2.04877e-19
c59 20 Vss 0.221837f
c60 17 Vss 0.180502f
c61 15 Vss 0.0247918f
c62 4 Vss 0.188411f
r63 93 98 0.441572
r64 92 94 0.655813
r65 92 93 9.04425
r66 88 98 0.174814
r67 84 98 0.441572
r68 52 94 3.33429
r69 47 88 3.33429
r70 40 57 1.16709
r71 40 84 22.1365
r72 40 44 0.0416786
r73 37 52 1.16709
r74 32 47 1.16709
r75 23 57 0.0476429
r76 21 23 0.326018
r77 21 23 0.1167
r78 20 24 0.652036
r79 20 23 6.7686
r80 17 57 0.357321
r81 15 23 0.326018
r82 15 17 0.40845
r83 8 37 0.123773
r84 6 32 0.123773
r85 4 24 5.1348
r86 2 17 4.72635
.ends

.subckt PM_G5_XOR3_N3_VSS 3 6 8 11 15 18 34 37 44 45 54 55 57 66 70 73 78 83 88
+ 93 98 107 112 121 123 124 125 130 131 136 142 145 154 155 156 Vss
c110 156 Vss 3.75522e-19
c111 155 Vss 3.91906e-19
c112 154 Vss 4.4306e-19
c113 142 Vss 0.00252991f
c114 136 Vss 0.00380695f
c115 131 Vss 8.45126e-19
c116 130 Vss 0.00638861f
c117 125 Vss 8.42189e-19
c118 124 Vss 0.0059194f
c119 123 Vss 0.00432257f
c120 121 Vss 0.00374747f
c121 112 Vss 0.00407665f
c122 107 Vss 0.00420294f
c123 98 Vss 0.00605485f
c124 93 Vss 0.00198064f
c125 88 Vss 8.56162e-19
c126 83 Vss 0.00102135f
c127 78 Vss 0.00266782f
c128 73 Vss 0.00352975f
c129 70 Vss 0.0100681f
c130 66 Vss 0.00715185f
c131 57 Vss 9.01088e-20
c132 55 Vss 0.0347733f
c133 54 Vss 0.0999406f
c134 45 Vss 0.035088f
c135 44 Vss 0.0994129f
c136 37 Vss 5.39995e-20
c137 35 Vss 0.0349058f
c138 34 Vss 0.100344f
c139 15 Vss 0.379408f
c140 11 Vss 0.379783f
c141 8 Vss 0.00143493f
c142 3 Vss 0.3841f
r143 143 156 0.494161
r144 143 145 6.62689
r145 142 150 0.652036
r146 142 145 0.833571
r147 138 156 0.128424
r148 137 155 0.494161
r149 136 146 0.652036
r150 136 137 7.46046
r151 132 155 0.128424
r152 130 156 0.494161
r153 130 131 15.8795
r154 126 154 0.0828784
r155 124 155 0.494161
r156 124 125 13.0037
r157 123 131 0.652036
r158 122 154 0.551426
r159 122 123 13.8373
r160 121 154 0.551426
r161 120 125 0.652036
r162 120 121 10.0029
r163 93 150 6.16843
r164 88 112 1.16709
r165 88 146 2.16729
r166 83 107 1.16709
r167 83 138 2.16729
r168 78 132 6.16843
r169 73 98 1.16709
r170 73 126 4.33978
r171 70 93 1.16709
r172 66 78 1.16709
r173 57 112 0.0476429
r174 55 57 1.45875
r175 54 58 0.652036
r176 54 57 1.45875
r177 51 55 0.652036
r178 47 107 0.0476429
r179 45 47 1.45875
r180 44 48 0.652036
r181 44 47 1.45875
r182 41 45 0.652036
r183 37 98 0.238214
r184 35 37 1.45875
r185 34 38 0.652036
r186 34 37 1.45875
r187 31 35 0.652036
r188 18 70 0.123773
r189 15 58 5.1348
r190 15 51 5.1348
r191 11 48 5.1348
r192 11 41 5.1348
r193 8 66 0.123773
r194 6 66 0.123773
r195 3 38 5.1348
r196 3 31 5.1348
.ends

.subckt PM_G5_XOR3_N3_CI 2 4 6 8 23 26 31 34 39 44 79 80 82 84 89 Vss
c52 95 Vss 8.92453e-20
c53 89 Vss 0.00607467f
c54 84 Vss 1.6915e-19
c55 83 Vss 1.82188e-19
c56 82 Vss 0.00167496f
c57 80 Vss 4.34795e-19
c58 79 Vss 0.00544906f
c59 44 Vss 7.72828e-19
c60 39 Vss 9.91594e-19
c61 34 Vss 0.00323815f
c62 31 Vss 0.00967911f
c63 26 Vss 0.00811165f
c64 23 Vss 0.00522928f
c65 4 Vss 0.00143493f
r66 90 95 0.494161
r67 89 91 0.652036
r68 89 90 10.3363
r69 85 95 0.128424
r70 83 95 0.494161
r71 83 84 1.50043
r72 82 84 0.652036
r73 81 82 6.46018
r74 79 81 0.652036
r75 79 80 19.1721
r76 75 80 0.652036
r77 44 91 3.41764
r78 39 85 3.41764
r79 34 75 8.62746
r80 31 44 1.16709
r81 26 39 1.16709
r82 23 34 1.16709
r83 8 31 0.123773
r84 6 26 0.123773
r85 4 23 0.123773
r86 2 23 0.123773
.ends

.subckt PM_G5_XOR3_N3_A 2 4 7 11 24 44 45 49 51 54 55 57 59 62 67 72 Vss
c67 72 Vss 0.00561856f
c68 67 Vss 0.00509443f
c69 59 Vss 9.40202e-19
c70 57 Vss 0.00665603f
c71 55 Vss 6.2663e-19
c72 54 Vss 0.00565582f
c73 51 Vss 0.00800572f
c74 49 Vss 0.135088f
c75 45 Vss 0.128114f
c76 44 Vss 1.14131e-19
c77 24 Vss 0.221923f
c78 21 Vss 0.18375f
c79 19 Vss 0.0247918f
c80 7 Vss 1.43819f
c81 4 Vss 0.194116f
r82 64 67 1.16709
r83 62 64 0.0416786
r84 59 62 0.833571
r85 57 72 1.16709
r86 55 57 9.66422
r87 53 55 0.655813
r88 53 54 10.4613
r89 52 59 0.0685365
r90 51 54 0.652036
r91 51 52 10.2113
r92 47 49 4.53833
r93 44 72 0.0238214
r94 44 45 2.26917
r95 41 44 2.26917
r96 36 49 0.00605528
r97 35 45 0.00605528
r98 32 47 0.00605528
r99 31 41 0.00605528
r100 27 67 0.0952857
r101 25 27 0.326018
r102 25 27 0.1167
r103 24 28 0.652036
r104 24 27 6.7686
r105 21 27 0.3335
r106 19 27 0.326018
r107 19 21 0.2334
r108 11 36 5.1348
r109 11 32 5.1348
r110 7 11 17.9718
r111 7 35 5.1348
r112 7 11 17.9718
r113 7 31 5.1348
r114 4 28 5.1348
r115 2 21 4.9014
.ends

.subckt PM_G5_XOR3_N3_BI 2 4 6 8 18 21 29 32 37 42 51 56 65 71 72 80 Vss
c62 80 Vss 3.85169e-19
c63 72 Vss 3.10144e-19
c64 71 Vss 7.91966e-19
c65 65 Vss 0.00115548f
c66 56 Vss 0.00255458f
c67 51 Vss 0.0023957f
c68 42 Vss 0.00128972f
c69 37 Vss 0.00247226f
c70 32 Vss 0.00178645f
c71 29 Vss 0.00520864f
c72 21 Vss 0.166484f
c73 6 Vss 0.166668f
c74 4 Vss 0.00143493f
r75 76 80 0.655813
r76 71 72 0.655813
r77 70 71 3.501
r78 65 70 0.655813
r79 42 56 1.16709
r80 42 72 2.00578
r81 37 51 1.16709
r82 37 80 12.0712
r83 37 65 2.00578
r84 32 76 3.33429
r85 29 32 1.16709
r86 21 56 0.50025
r87 18 51 0.50025
r88 8 21 4.37625
r89 6 18 4.37625
r90 4 29 0.123773
r91 2 29 0.123773
.ends

.subckt PM_G5_XOR3_N3_AI 2 4 7 11 31 37 43 46 51 60 73 79 Vss
c44 79 Vss 2.91008e-19
c45 73 Vss 0.00515518f
c46 60 Vss 0.0064096f
c47 51 Vss 0.00263851f
c48 46 Vss 0.0021137f
c49 43 Vss 0.0046119f
c50 37 Vss 0.12791f
c51 31 Vss 0.131715f
c52 7 Vss 1.42572f
c53 4 Vss 0.00143493f
r54 75 79 0.652036
r55 73 79 13.7539
r56 51 60 1.16709
r57 51 73 2.75079
r58 46 75 6.16843
r59 43 46 1.16709
r60 36 60 0.0238214
r61 36 37 2.334
r62 33 36 2.20433
r63 29 31 4.53833
r64 26 37 0.00605528
r65 25 31 0.00605528
r66 22 33 0.00605528
r67 21 29 0.00605528
r68 11 26 5.1348
r69 11 22 5.1348
r70 7 11 17.9718
r71 7 25 5.1348
r72 7 11 17.9718
r73 7 21 5.1348
r74 4 43 0.123773
r75 2 43 0.123773
.ends

.subckt PM_G5_XOR3_N3_B 2 4 6 8 16 17 24 26 33 38 42 45 50 55 60 65 73 74 80 86
+ 91 92 Vss
c69 92 Vss 2.0377e-19
c70 91 Vss 6.9543e-19
c71 86 Vss 8.47373e-19
c72 80 Vss 9.51093e-19
c73 74 Vss 5.10711e-19
c74 73 Vss 0.00481884f
c75 65 Vss 0.00266055f
c76 60 Vss 0.00231285f
c77 55 Vss 0.00437951f
c78 50 Vss 0.00146415f
c79 45 Vss 4.84439e-19
c80 42 Vss 7.72719e-19
c81 38 Vss 7.58106e-19
c82 33 Vss 9.01088e-20
c83 26 Vss 0.166484f
c84 24 Vss 1.01938e-19
c85 20 Vss 0.0247918f
c86 17 Vss 0.0340157f
c87 16 Vss 0.186033f
c88 8 Vss 0.166484f
c89 4 Vss 0.180512f
c90 2 Vss 0.191454f
r91 90 92 0.655813
r92 90 91 3.501
r93 86 91 0.655813
r94 73 80 0.0685365
r95 73 74 10.3363
r96 69 74 0.652036
r97 50 65 1.16709
r98 50 92 2.00578
r99 45 60 1.16709
r100 45 86 2.00578
r101 45 80 2.04225
r102 38 55 1.16709
r103 38 69 2.20896
r104 38 42 0.0729375
r105 36 55 0.0476429
r106 33 65 0.50025
r107 26 60 0.50025
r108 24 55 0.357321
r109 20 36 0.326018
r110 20 24 0.40845
r111 17 36 6.7686
r112 16 36 0.326018
r113 16 36 0.1167
r114 13 17 0.652036
r115 8 33 4.37625
r116 6 26 4.37625
r117 4 24 4.72635
r118 2 13 5.1348
.ends

.subckt PM_G5_XOR3_N3_Z 2 4 6 8 23 27 30 33 Vss
c32 30 Vss 0.00377706f
c33 27 Vss 0.00795274f
c34 23 Vss 0.00720799f
c35 8 Vss 0.00143493f
c36 6 Vss 0.00334888f
r37 33 35 7.21039
r38 30 40 1.16709
r39 30 33 5.62661
r40 27 35 1.16709
r41 23 40 0.05
r42 8 27 0.123773
r43 6 23 0.123773
r44 4 27 0.123773
r45 2 23 0.123773
.ends

.subckt G5_XOR3_N3  VDD C VSS A B Z
*
* Z	Z
* B	B
* A	A
* VSS	VSS
* C	C
* VDD	VDD
XI25.X0 N_CI_XI25.X0_D N_VSS_XI25.X0_PGD N_C_XI25.X0_CG N_VSS_XI25.X0_PGD
+ N_VDD_XI25.X0_S TIGFET_HPNW12
XI22.X0 N_CI_XI22.X0_D N_VDD_XI22.X0_PGD N_C_XI22.X0_CG N_VDD_XI22.X0_PGD
+ N_VSS_XI22.X0_S TIGFET_HPNW12
XI21.X0 N_BI_XI21.X0_D N_VDD_XI21.X0_PGD N_B_XI21.X0_CG N_VDD_XI21.X0_PGD
+ N_VSS_XI21.X0_S TIGFET_HPNW12
XI23.X0 N_AI_XI23.X0_D N_VSS_XI23.X0_PGD N_A_XI23.X0_CG N_VSS_XI23.X0_PGD
+ N_VDD_XI23.X0_S TIGFET_HPNW12
XI24.X0 N_BI_XI24.X0_D N_VSS_XI24.X0_PGD N_B_XI24.X0_CG N_VSS_XI24.X0_PGD
+ N_VDD_XI24.X0_S TIGFET_HPNW12
XI20.X0 N_AI_XI20.X0_D N_VDD_XI20.X0_PGD N_A_XI20.X0_CG N_VDD_XI20.X0_PGD
+ N_VSS_XI20.X0_S TIGFET_HPNW12
XI29.X0 N_Z_XI29.X0_D N_AI_XI29.X0_PGD N_BI_XI29.X0_CG N_AI_XI29.X0_PGD
+ N_C_XI29.X0_S TIGFET_HPNW12
XI27.X0 N_Z_XI27.X0_D N_AI_XI27.X0_PGD N_B_XI27.X0_CG N_AI_XI27.X0_PGD
+ N_CI_XI27.X0_S TIGFET_HPNW12
XI28.X0 N_Z_XI28.X0_D N_A_XI28.X0_PGD N_B_XI28.X0_CG N_A_XI28.X0_PGD
+ N_C_XI28.X0_S TIGFET_HPNW12
XI26.X0 N_Z_XI26.X0_D N_A_XI26.X0_PGD N_BI_XI26.X0_CG N_A_XI26.X0_PGD
+ N_CI_XI26.X0_S TIGFET_HPNW12
*
x_PM_G5_XOR3_N3_VDD N_VDD_XI25.X0_S N_VDD_XI22.X0_PGD N_VDD_XI21.X0_PGD
+ N_VDD_XI23.X0_S N_VDD_XI24.X0_S N_VDD_XI20.X0_PGD N_VDD_c_111_p N_VDD_c_19_p
+ N_VDD_c_24_p N_VDD_c_4_p N_VDD_c_100_p N_VDD_c_20_p N_VDD_c_74_p N_VDD_c_101_p
+ N_VDD_c_6_p N_VDD_c_7_p N_VDD_c_13_p N_VDD_c_5_p N_VDD_c_61_p N_VDD_c_29_p
+ N_VDD_c_62_p N_VDD_c_30_p N_VDD_c_16_p N_VDD_c_63_p N_VDD_c_21_p N_VDD_c_10_p
+ N_VDD_c_25_p N_VDD_c_37_p N_VDD_c_11_p N_VDD_c_57_p VDD N_VDD_c_65_p
+ N_VDD_c_69_p N_VDD_c_2_p N_VDD_c_42_p N_VDD_c_38_p Vss PM_G5_XOR3_N3_VDD
x_PM_G5_XOR3_N3_C N_C_XI25.X0_CG N_C_XI22.X0_CG N_C_XI29.X0_S N_C_XI28.X0_S
+ N_C_c_130_p N_C_c_116_n N_C_c_126_p N_C_c_119_n N_C_c_157_p N_C_c_120_n C
+ N_C_c_127_p N_C_c_159_p N_C_c_122_n N_C_c_123_n N_C_c_145_p N_C_c_146_p Vss
+ PM_G5_XOR3_N3_C
x_PM_G5_XOR3_N3_VSS N_VSS_XI25.X0_PGD N_VSS_XI22.X0_S N_VSS_XI21.X0_S
+ N_VSS_XI23.X0_PGD N_VSS_XI24.X0_PGD N_VSS_XI20.X0_S N_VSS_c_170_n
+ N_VSS_c_226_n N_VSS_c_171_n N_VSS_c_173_n N_VSS_c_174_n N_VSS_c_175_n
+ N_VSS_c_269_p N_VSS_c_177_n N_VSS_c_238_p N_VSS_c_178_n N_VSS_c_183_n
+ N_VSS_c_186_n N_VSS_c_190_n N_VSS_c_194_n N_VSS_c_195_n N_VSS_c_198_n
+ N_VSS_c_202_n N_VSS_c_206_n N_VSS_c_209_n N_VSS_c_211_n N_VSS_c_212_n
+ N_VSS_c_213_n N_VSS_c_217_n N_VSS_c_218_n N_VSS_c_221_n VSS N_VSS_c_222_n
+ N_VSS_c_223_n N_VSS_c_224_n Vss PM_G5_XOR3_N3_VSS
x_PM_G5_XOR3_N3_CI N_CI_XI25.X0_D N_CI_XI22.X0_D N_CI_XI27.X0_S N_CI_XI26.X0_S
+ N_CI_c_273_n N_CI_c_286_n N_CI_c_317_p N_CI_c_275_n N_CI_c_292_n N_CI_c_319_p
+ N_CI_c_279_n N_CI_c_295_n N_CI_c_296_n N_CI_c_308_p N_CI_c_302_p Vss
+ PM_G5_XOR3_N3_CI
x_PM_G5_XOR3_N3_A N_A_XI23.X0_CG N_A_XI20.X0_CG N_A_XI28.X0_PGD N_A_XI26.X0_PGD
+ N_A_c_325_n N_A_c_374_p N_A_c_365_p N_A_c_367_p N_A_c_326_n N_A_c_332_n
+ N_A_c_333_n N_A_c_340_n N_A_c_334_n A N_A_c_335_n N_A_c_378_p Vss
+ PM_G5_XOR3_N3_A
x_PM_G5_XOR3_N3_BI N_BI_XI21.X0_D N_BI_XI24.X0_D N_BI_XI29.X0_CG N_BI_XI26.X0_CG
+ N_BI_c_412_n N_BI_c_413_n N_BI_c_392_n N_BI_c_395_n N_BI_c_399_n N_BI_c_410_n
+ N_BI_c_418_n N_BI_c_419_n N_BI_c_402_n N_BI_c_440_p N_BI_c_428_p N_BI_c_403_n
+ Vss PM_G5_XOR3_N3_BI
x_PM_G5_XOR3_N3_AI N_AI_XI23.X0_D N_AI_XI20.X0_D N_AI_XI29.X0_PGD
+ N_AI_XI27.X0_PGD N_AI_c_465_n N_AI_c_455_n N_AI_c_456_n N_AI_c_458_n
+ N_AI_c_471_n N_AI_c_492_p N_AI_c_463_n N_AI_c_473_n Vss PM_G5_XOR3_N3_AI
x_PM_G5_XOR3_N3_B N_B_XI21.X0_CG N_B_XI24.X0_CG N_B_XI27.X0_CG N_B_XI28.X0_CG
+ N_B_c_499_n N_B_c_500_n N_B_c_507_n N_B_c_557_n N_B_c_521_n N_B_c_501_n B
+ N_B_c_537_n N_B_c_512_n N_B_c_509_n N_B_c_541_n N_B_c_529_n N_B_c_502_n
+ N_B_c_514_n N_B_c_548_n N_B_c_504_n N_B_c_554_n N_B_c_505_n Vss
+ PM_G5_XOR3_N3_B
x_PM_G5_XOR3_N3_Z N_Z_XI29.X0_D N_Z_XI27.X0_D N_Z_XI28.X0_D N_Z_XI26.X0_D
+ N_Z_c_567_n N_Z_c_574_n N_Z_c_571_n Z Vss PM_G5_XOR3_N3_Z
cc_1 N_VDD_XI21.X0_PGD N_C_XI22.X0_CG 0.00111653f
cc_2 N_VDD_c_2_p N_C_XI22.X0_CG 0.00108697f
cc_3 N_VDD_XI22.X0_PGD N_C_c_116_n 4.20258e-19
cc_4 N_VDD_c_4_p N_C_c_116_n 0.00111653f
cc_5 N_VDD_c_5_p N_C_c_116_n 0.00135138f
cc_6 N_VDD_c_6_p N_C_c_119_n 3.43419e-19
cc_7 N_VDD_c_7_p N_C_c_120_n 4.76491e-19
cc_8 N_VDD_c_5_p N_C_c_120_n 0.00161703f
cc_9 N_VDD_c_5_p N_C_c_122_n 2.84771e-19
cc_10 N_VDD_c_10_p N_C_c_123_n 5.24769e-19
cc_11 N_VDD_c_11_p N_C_c_123_n 8.43519e-19
cc_12 N_VDD_XI22.X0_PGD N_VSS_XI25.X0_PGD 0.00200994f
cc_13 N_VDD_c_13_p N_VSS_XI25.X0_PGD 4.18763e-19
cc_14 N_VDD_XI21.X0_PGD N_VSS_XI23.X0_PGD 2.44446e-19
cc_15 N_VDD_XI20.X0_PGD N_VSS_XI23.X0_PGD 0.00201012f
cc_16 N_VDD_c_16_p N_VSS_XI23.X0_PGD 4.21402e-19
cc_17 N_VDD_XI21.X0_PGD N_VSS_XI24.X0_PGD 0.00200584f
cc_18 N_VDD_XI20.X0_PGD N_VSS_XI24.X0_PGD 2.31301e-19
cc_19 N_VDD_c_19_p N_VSS_c_170_n 0.00200994f
cc_20 N_VDD_c_20_p N_VSS_c_171_n 0.00201012f
cc_21 N_VDD_c_21_p N_VSS_c_171_n 3.00545e-19
cc_22 N_VDD_c_21_p N_VSS_c_173_n 3.89167e-19
cc_23 N_VDD_c_11_p N_VSS_c_174_n 2.35465e-19
cc_24 N_VDD_c_24_p N_VSS_c_175_n 0.00200584f
cc_25 N_VDD_c_25_p N_VSS_c_175_n 3.89167e-19
cc_26 N_VDD_c_5_p N_VSS_c_177_n 2.74986e-19
cc_27 N_VDD_c_13_p N_VSS_c_178_n 4.32468e-19
cc_28 N_VDD_c_5_p N_VSS_c_178_n 3.08724e-19
cc_29 N_VDD_c_29_p N_VSS_c_178_n 0.00111881f
cc_30 N_VDD_c_30_p N_VSS_c_178_n 3.98949e-19
cc_31 N_VDD_c_2_p N_VSS_c_178_n 3.48267e-19
cc_32 N_VDD_c_5_p N_VSS_c_183_n 2.9533e-19
cc_33 N_VDD_c_10_p N_VSS_c_183_n 7.43603e-19
cc_34 N_VDD_c_11_p N_VSS_c_183_n 8.20353e-19
cc_35 N_VDD_c_16_p N_VSS_c_186_n 6.74818e-19
cc_36 N_VDD_c_21_p N_VSS_c_186_n 0.00161703f
cc_37 N_VDD_c_37_p N_VSS_c_186_n 8.6926e-19
cc_38 N_VDD_c_38_p N_VSS_c_186_n 3.48267e-19
cc_39 N_VDD_c_10_p N_VSS_c_190_n 6.78479e-19
cc_40 N_VDD_c_25_p N_VSS_c_190_n 0.00161703f
cc_41 N_VDD_c_11_p N_VSS_c_190_n 0.0024227f
cc_42 N_VDD_c_42_p N_VSS_c_190_n 3.48267e-19
cc_43 N_VDD_c_37_p N_VSS_c_194_n 7.32365e-19
cc_44 N_VDD_c_13_p N_VSS_c_195_n 4.41003e-19
cc_45 N_VDD_c_30_p N_VSS_c_195_n 3.89161e-19
cc_46 N_VDD_c_2_p N_VSS_c_195_n 7.99831e-19
cc_47 N_VDD_c_16_p N_VSS_c_198_n 3.48267e-19
cc_48 N_VDD_c_21_p N_VSS_c_198_n 2.26455e-19
cc_49 N_VDD_c_37_p N_VSS_c_198_n 3.99794e-19
cc_50 N_VDD_c_38_p N_VSS_c_198_n 6.489e-19
cc_51 N_VDD_c_10_p N_VSS_c_202_n 3.82294e-19
cc_52 N_VDD_c_25_p N_VSS_c_202_n 2.26455e-19
cc_53 N_VDD_c_11_p N_VSS_c_202_n 9.55109e-19
cc_54 N_VDD_c_42_p N_VSS_c_202_n 6.46219e-19
cc_55 N_VDD_c_7_p N_VSS_c_206_n 0.00419405f
cc_56 N_VDD_c_13_p N_VSS_c_206_n 0.00330716f
cc_57 N_VDD_c_57_p N_VSS_c_206_n 0.0010705f
cc_58 N_VDD_c_13_p N_VSS_c_209_n 0.00977753f
cc_59 N_VDD_c_30_p N_VSS_c_209_n 0.00139461f
cc_60 N_VDD_c_5_p N_VSS_c_211_n 0.0097003f
cc_61 N_VDD_c_61_p N_VSS_c_212_n 0.00107633f
cc_62 N_VDD_c_62_p N_VSS_c_213_n 0.00839359f
cc_63 N_VDD_c_63_p N_VSS_c_213_n 6.54257e-19
cc_64 N_VDD_c_21_p N_VSS_c_213_n 0.00374326f
cc_65 N_VDD_c_65_p N_VSS_c_213_n 0.00149946f
cc_66 N_VDD_c_13_p N_VSS_c_217_n 0.00107845f
cc_67 N_VDD_c_5_p N_VSS_c_218_n 0.00143483f
cc_68 N_VDD_c_25_p N_VSS_c_218_n 0.00612925f
cc_69 N_VDD_c_69_p N_VSS_c_218_n 9.53204e-19
cc_70 N_VDD_c_21_p N_VSS_c_221_n 0.00550311f
cc_71 N_VDD_c_13_p N_VSS_c_222_n 0.00112682f
cc_72 N_VDD_c_5_p N_VSS_c_223_n 0.00111918f
cc_73 N_VDD_c_21_p N_VSS_c_224_n 7.74609e-19
cc_74 N_VDD_c_74_p N_CI_c_273_n 3.43419e-19
cc_75 N_VDD_c_29_p N_CI_c_273_n 3.72199e-19
cc_76 N_VDD_c_74_p N_CI_c_275_n 3.48267e-19
cc_77 N_VDD_c_5_p N_CI_c_275_n 3.21336e-19
cc_78 N_VDD_c_29_p N_CI_c_275_n 5.226e-19
cc_79 N_VDD_c_30_p N_CI_c_275_n 0.00102111f
cc_80 N_VDD_c_30_p N_CI_c_279_n 7.25102e-19
cc_81 N_VDD_c_63_p N_CI_c_279_n 7.87445e-19
cc_82 N_VDD_XI20.X0_PGD N_A_c_325_n 3.97033e-19
cc_83 N_VDD_XI20.X0_PGD N_A_c_326_n 2.7861e-19
cc_84 N_VDD_c_6_p N_A_c_326_n 2.23042e-19
cc_85 N_VDD_c_21_p N_A_c_326_n 3.21337e-19
cc_86 N_VDD_c_37_p N_A_c_326_n 2.93421e-19
cc_87 N_VDD_c_11_p N_A_c_326_n 3.31604e-19
cc_88 N_VDD_c_38_p N_A_c_326_n 2.04325e-19
cc_89 N_VDD_c_6_p N_A_c_332_n 9.18655e-19
cc_90 N_VDD_c_11_p N_A_c_333_n 0.00704792f
cc_91 N_VDD_c_30_p N_A_c_334_n 0.00104803f
cc_92 N_VDD_c_30_p N_A_c_335_n 5.71346e-19
cc_93 N_VDD_c_6_p N_BI_c_392_n 3.43419e-19
cc_94 N_VDD_c_25_p N_BI_c_392_n 2.74986e-19
cc_95 N_VDD_c_11_p N_BI_c_392_n 3.48267e-19
cc_96 N_VDD_c_6_p N_BI_c_395_n 3.48267e-19
cc_97 N_VDD_c_25_p N_BI_c_395_n 2.9533e-19
cc_98 N_VDD_c_11_p N_BI_c_395_n 4.99861e-19
cc_99 N_VDD_XI20.X0_PGD N_AI_XI29.X0_PGD 3.2392e-19
cc_100 N_VDD_c_100_p N_AI_c_455_n 3.2392e-19
cc_101 N_VDD_c_101_p N_AI_c_456_n 3.43419e-19
cc_102 N_VDD_c_63_p N_AI_c_456_n 3.73302e-19
cc_103 N_VDD_c_101_p N_AI_c_458_n 3.48267e-19
cc_104 N_VDD_c_16_p N_AI_c_458_n 3.24512e-19
cc_105 N_VDD_c_63_p N_AI_c_458_n 5.23123e-19
cc_106 N_VDD_c_21_p N_AI_c_458_n 3.21336e-19
cc_107 N_VDD_c_37_p N_AI_c_458_n 5.55696e-19
cc_108 N_VDD_c_21_p N_AI_c_463_n 4.73141e-19
cc_109 N_VDD_XI22.X0_PGD N_B_XI21.X0_CG 0.00111821f
cc_110 N_VDD_XI21.X0_PGD N_B_c_499_n 4.01531e-19
cc_111 N_VDD_c_111_p N_B_c_500_n 0.00111821f
cc_112 N_VDD_c_30_p N_B_c_501_n 7.28643e-19
cc_113 N_VDD_c_11_p N_B_c_502_n 2.93412e-19
cc_114 N_C_c_116_n N_VSS_XI25.X0_PGD 4.20258e-19
cc_115 N_C_c_126_p N_VSS_c_226_n 2.76939e-19
cc_116 N_C_c_127_p N_VSS_c_183_n 7.31268e-19
cc_117 N_C_c_123_n N_VSS_c_183_n 0.00201674f
cc_118 N_C_c_123_n N_VSS_c_190_n 0.00162673f
cc_119 N_C_c_130_p N_VSS_c_195_n 0.0041528f
cc_120 N_C_c_120_n N_VSS_c_206_n 4.01014e-19
cc_121 N_C_c_123_n N_VSS_c_206_n 2.67373e-19
cc_122 N_C_c_120_n N_VSS_c_211_n 0.00171716f
cc_123 N_C_c_123_n N_VSS_c_211_n 0.00318423f
cc_124 N_C_c_123_n N_VSS_c_218_n 0.00194657f
cc_125 N_C_c_116_n N_CI_c_273_n 7.69306e-19
cc_126 N_C_c_123_n N_CI_c_275_n 7.41148e-19
cc_127 N_C_c_123_n N_CI_c_279_n 0.00247018f
cc_128 N_C_c_123_n N_A_c_326_n 2.96232e-19
cc_129 N_C_c_119_n N_A_c_332_n 8.20481e-19
cc_130 N_C_c_127_p N_A_c_332_n 0.00202163f
cc_131 N_C_c_123_n N_A_c_333_n 5.81147e-19
cc_132 N_C_c_127_p N_A_c_340_n 0.00128177f
cc_133 N_C_c_123_n N_A_c_340_n 4.89987e-19
cc_134 N_C_c_145_p N_A_c_340_n 0.00290875f
cc_135 N_C_c_146_p N_A_c_340_n 3.99251e-19
cc_136 N_C_c_123_n N_BI_c_395_n 7.95957e-19
cc_137 N_C_c_127_p N_BI_c_399_n 8.44326e-19
cc_138 N_C_c_123_n N_BI_c_399_n 0.00305118f
cc_139 N_C_c_145_p N_BI_c_399_n 4.85495e-19
cc_140 N_C_c_145_p N_BI_c_402_n 7.42134e-19
cc_141 N_C_c_123_n N_BI_c_403_n 5.13569e-19
cc_142 N_C_c_127_p N_B_c_502_n 6.36664e-19
cc_143 N_C_c_145_p N_B_c_504_n 3.34841e-19
cc_144 N_C_c_145_p N_B_c_505_n 0.0012842f
cc_145 N_C_c_119_n N_Z_c_567_n 3.43419e-19
cc_146 N_C_c_157_p N_Z_c_567_n 3.43419e-19
cc_147 N_C_c_127_p N_Z_c_567_n 3.48267e-19
cc_148 N_C_c_159_p N_Z_c_567_n 3.48267e-19
cc_149 N_C_c_157_p N_Z_c_571_n 3.48267e-19
cc_150 N_C_c_127_p N_Z_c_571_n 6.09821e-19
cc_151 N_C_c_159_p N_Z_c_571_n 5.71987e-19
cc_152 N_VSS_c_177_n N_CI_c_273_n 3.43419e-19
cc_153 N_VSS_c_183_n N_CI_c_273_n 3.48267e-19
cc_154 N_VSS_c_238_p N_CI_c_286_n 3.43419e-19
cc_155 N_VSS_c_177_n N_CI_c_275_n 3.48267e-19
cc_156 N_VSS_c_178_n N_CI_c_275_n 5.88914e-19
cc_157 N_VSS_c_183_n N_CI_c_275_n 8.10527e-19
cc_158 N_VSS_c_206_n N_CI_c_275_n 7.39772e-19
cc_159 N_VSS_c_209_n N_CI_c_275_n 9.66332e-19
cc_160 N_VSS_c_194_n N_CI_c_292_n 8.792e-19
cc_161 N_VSS_c_186_n N_CI_c_279_n 3.71583e-19
cc_162 N_VSS_c_221_n N_CI_c_279_n 4.92938e-19
cc_163 N_VSS_c_213_n N_CI_c_295_n 0.00161605f
cc_164 N_VSS_c_194_n N_CI_c_296_n 0.00179737f
cc_165 N_VSS_XI23.X0_PGD N_A_c_325_n 3.97033e-19
cc_166 N_VSS_c_194_n N_A_c_326_n 6.39942e-19
cc_167 N_VSS_c_221_n N_A_c_326_n 3.79499e-19
cc_168 N_VSS_c_198_n N_A_c_334_n 2.09367e-19
cc_169 N_VSS_c_186_n N_A_c_335_n 2.04211e-19
cc_170 N_VSS_c_198_n N_A_c_335_n 4.89964e-19
cc_171 N_VSS_c_177_n N_BI_c_392_n 3.43419e-19
cc_172 N_VSS_c_177_n N_BI_c_395_n 3.48267e-19
cc_173 N_VSS_c_183_n N_BI_c_395_n 8.48361e-19
cc_174 N_VSS_XI24.X0_PGD N_AI_XI29.X0_PGD 2.79882e-19
cc_175 N_VSS_c_174_n N_AI_c_465_n 2.79882e-19
cc_176 N_VSS_c_238_p N_AI_c_456_n 3.43419e-19
cc_177 N_VSS_c_238_p N_AI_c_458_n 3.48267e-19
cc_178 N_VSS_c_186_n N_AI_c_458_n 0.00108072f
cc_179 N_VSS_c_194_n N_AI_c_458_n 0.00227024f
cc_180 N_VSS_c_209_n N_AI_c_458_n 7.83107e-19
cc_181 N_VSS_c_194_n N_AI_c_471_n 0.00125351f
cc_182 N_VSS_c_221_n N_AI_c_463_n 0.00560835f
cc_183 N_VSS_c_221_n N_AI_c_473_n 0.00192498f
cc_184 N_VSS_XI24.X0_PGD N_B_c_499_n 4.01531e-19
cc_185 N_VSS_c_269_p N_B_c_507_n 5.35095e-19
cc_186 N_VSS_c_202_n B 2.15082e-19
cc_187 N_VSS_c_190_n N_B_c_509_n 2.15082e-19
cc_188 N_VSS_c_194_n N_B_c_502_n 2.6453e-19
cc_189 N_CI_c_279_n N_A_c_326_n 0.00190043f
cc_190 N_CI_c_279_n N_A_c_334_n 3.93937e-19
cc_191 N_CI_c_275_n N_BI_c_395_n 0.00116552f
cc_192 N_CI_c_292_n N_BI_c_399_n 2.45753e-19
cc_193 N_CI_c_279_n N_BI_c_399_n 0.00333331f
cc_194 N_CI_c_302_p N_BI_c_410_n 7.0273e-19
cc_195 N_CI_c_279_n N_BI_c_403_n 0.00154189f
cc_196 N_CI_c_279_n N_AI_c_458_n 9.328e-19
cc_197 N_CI_c_296_n N_AI_c_458_n 0.00145606f
cc_198 N_CI_c_302_p N_AI_c_471_n 0.00147513f
cc_199 N_CI_c_279_n N_AI_c_463_n 0.00163581f
cc_200 N_CI_c_308_p N_AI_c_463_n 0.00486757f
cc_201 N_CI_c_302_p N_AI_c_463_n 0.00259545f
cc_202 N_CI_c_275_n N_B_c_501_n 5.60809e-19
cc_203 N_CI_c_302_p N_B_c_512_n 5.08667e-19
cc_204 N_CI_c_292_n N_B_c_502_n 7.44351e-19
cc_205 N_CI_c_279_n N_B_c_514_n 0.00125143f
cc_206 N_CI_c_279_n N_B_c_504_n 4.54745e-19
cc_207 N_CI_c_302_p N_B_c_504_n 0.00126146f
cc_208 N_CI_c_286_n N_Z_c_574_n 3.43419e-19
cc_209 N_CI_c_317_p N_Z_c_574_n 3.43419e-19
cc_210 N_CI_c_292_n N_Z_c_574_n 3.48267e-19
cc_211 N_CI_c_319_p N_Z_c_574_n 3.48267e-19
cc_212 N_CI_c_286_n N_Z_c_571_n 3.48267e-19
cc_213 N_CI_c_317_p N_Z_c_571_n 3.48267e-19
cc_214 N_CI_c_292_n N_Z_c_571_n 5.71987e-19
cc_215 N_CI_c_319_p N_Z_c_571_n 5.71987e-19
cc_216 N_CI_c_279_n N_Z_c_571_n 6.3795e-19
cc_217 N_A_c_340_n N_BI_c_412_n 2.09474e-19
cc_218 N_A_XI28.X0_PGD N_BI_c_413_n 9.65637e-19
cc_219 N_A_c_326_n N_BI_c_395_n 3.45209e-19
cc_220 N_A_c_332_n N_BI_c_395_n 6.2874e-19
cc_221 N_A_c_332_n N_BI_c_399_n 0.00115936f
cc_222 N_A_c_340_n N_BI_c_399_n 6.34965e-19
cc_223 N_A_c_332_n N_BI_c_418_n 3.37713e-19
cc_224 N_A_XI28.X0_PGD N_BI_c_419_n 0.00133285f
cc_225 N_A_c_340_n N_BI_c_402_n 7.80641e-19
cc_226 N_A_c_326_n N_BI_c_403_n 4.18438e-19
cc_227 N_A_XI28.X0_PGD N_AI_XI29.X0_PGD 0.0174159f
cc_228 N_A_c_332_n N_AI_XI29.X0_PGD 9.45724e-19
cc_229 N_A_c_340_n N_AI_XI29.X0_PGD 7.67512e-19
cc_230 N_A_c_365_p N_AI_c_465_n 0.00199603f
cc_231 N_A_c_340_n N_AI_c_465_n 0.00129811f
cc_232 N_A_c_367_p N_AI_c_455_n 0.00201004f
cc_233 N_A_c_325_n N_AI_c_456_n 6.90199e-19
cc_234 N_A_c_326_n N_AI_c_458_n 5.93425e-19
cc_235 N_A_XI28.X0_PGD N_B_XI28.X0_CG 9.65637e-19
cc_236 N_A_c_325_n N_B_c_499_n 0.00358744f
cc_237 N_A_c_326_n N_B_c_499_n 8.32052e-19
cc_238 N_A_c_335_n N_B_c_500_n 7.41063e-19
cc_239 N_A_c_374_p N_B_c_521_n 5.35095e-19
cc_240 N_A_c_332_n N_B_c_501_n 6.26711e-19
cc_241 N_A_c_326_n B 8.224e-19
cc_242 N_A_c_332_n B 5.04818e-19
cc_243 N_A_c_378_p N_B_c_512_n 2.15082e-19
cc_244 N_A_c_325_n N_B_c_509_n 0.00108715f
cc_245 N_A_c_326_n N_B_c_509_n 6.90512e-19
cc_246 N_A_c_332_n N_B_c_509_n 6.85754e-19
cc_247 N_A_XI28.X0_PGD N_B_c_529_n 0.00133285f
cc_248 N_A_c_340_n N_B_c_529_n 2.15082e-19
cc_249 N_A_c_326_n N_B_c_502_n 0.00340226f
cc_250 N_A_c_332_n N_B_c_502_n 0.00192865f
cc_251 N_A_c_340_n N_B_c_502_n 6.44056e-19
cc_252 N_A_c_326_n N_B_c_514_n 5.44597e-19
cc_253 N_A_c_340_n N_Z_c_567_n 5.87699e-19
cc_254 N_A_XI28.X0_PGD N_Z_c_571_n 7.94638e-19
cc_255 N_A_c_332_n N_Z_c_571_n 0.00175701f
cc_256 N_A_c_340_n N_Z_c_571_n 0.00103031f
cc_257 N_BI_XI29.X0_CG N_AI_XI29.X0_PGD 9.47088e-19
cc_258 N_BI_c_418_n N_AI_XI29.X0_PGD 0.00133285f
cc_259 N_BI_c_399_n N_AI_c_463_n 8.39468e-19
cc_260 N_BI_c_392_n N_B_c_499_n 6.90199e-19
cc_261 N_BI_c_399_n N_B_c_501_n 0.00133142f
cc_262 N_BI_c_399_n N_B_c_537_n 5.44238e-19
cc_263 N_BI_c_428_p N_B_c_537_n 3.08318e-19
cc_264 N_BI_c_410_n N_B_c_512_n 0.00187472f
cc_265 N_BI_c_402_n N_B_c_512_n 0.00165773f
cc_266 N_BI_c_399_n N_B_c_541_n 4.56568e-19
cc_267 N_BI_c_418_n N_B_c_541_n 0.00266356f
cc_268 N_BI_c_419_n N_B_c_541_n 7.16621e-19
cc_269 N_BI_c_410_n N_B_c_529_n 4.62769e-19
cc_270 N_BI_c_418_n N_B_c_529_n 6.17967e-19
cc_271 N_BI_c_419_n N_B_c_529_n 0.00243633f
cc_272 N_BI_c_399_n N_B_c_502_n 0.00398399f
cc_273 N_BI_c_399_n N_B_c_548_n 3.07174e-19
cc_274 N_BI_c_402_n N_B_c_548_n 0.00126004f
cc_275 N_BI_c_440_p N_B_c_548_n 0.00342237f
cc_276 N_BI_c_399_n N_B_c_504_n 5.09978e-19
cc_277 N_BI_c_402_n N_B_c_504_n 9.4756e-19
cc_278 N_BI_c_428_p N_B_c_504_n 8.92139e-19
cc_279 N_BI_c_440_p N_B_c_554_n 0.00210118f
cc_280 N_BI_c_399_n N_B_c_505_n 0.00143025f
cc_281 N_BI_c_402_n N_B_c_505_n 9.46104e-19
cc_282 N_BI_c_399_n N_Z_c_571_n 0.00138952f
cc_283 N_BI_c_410_n N_Z_c_571_n 0.00141294f
cc_284 N_BI_c_418_n N_Z_c_571_n 8.66889e-19
cc_285 N_BI_c_419_n N_Z_c_571_n 8.66889e-19
cc_286 N_BI_c_402_n N_Z_c_571_n 0.00105522f
cc_287 N_BI_c_440_p N_Z_c_571_n 0.00212989f
cc_288 N_BI_c_428_p N_Z_c_571_n 0.00104995f
cc_289 N_AI_XI29.X0_PGD N_B_c_557_n 9.65637e-19
cc_290 N_AI_c_492_p N_B_c_537_n 2.15082e-19
cc_291 N_AI_XI29.X0_PGD N_B_c_541_n 0.00133285f
cc_292 N_AI_c_471_n N_B_c_541_n 2.15082e-19
cc_293 N_AI_c_492_p N_B_c_541_n 5.05931e-19
cc_294 N_AI_c_463_n N_B_c_502_n 4.67711e-19
cc_295 N_AI_XI29.X0_PGD N_Z_c_571_n 4.32017e-19
cc_296 N_B_c_537_n N_Z_c_571_n 0.00157325f
cc_297 N_B_c_512_n N_Z_c_571_n 0.00138952f
cc_298 N_B_c_529_n N_Z_c_571_n 8.66889e-19
cc_299 N_B_c_548_n N_Z_c_571_n 4.69528e-19
*
.ends
*
*
.subckt XOR3_HPNW12 A B C Y VDD VSS
xgate (VDD C VSS A B Y) G5_XOR3_N3
.ends
